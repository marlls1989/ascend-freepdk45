
.SUBCKT FILLTIE VDD VSS
*.PININFO VDD:P VSS:G
.ENDS
******************************************************************************
*                                                                            *
* End of file.                                                               *
*                                                                            *
******************************************************************************

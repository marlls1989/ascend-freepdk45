
VERSION 5.6 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 

MACRO ACELEM1X1
  CLASS CORE ;
  FOREIGN ACELEM1X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.595 0.825 0.805 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.130 0.875 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.890 0.260 1.150 0.525 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038850 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.245 1.665 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.980 0.130 1.485 ;
        RECT 0.130 1.315 0.795 1.485 ;
        RECT 0.795 1.290 0.930 1.485 ;
        RECT 0.930 1.315 1.395 1.485 ;
        RECT 1.395 0.950 1.485 1.485 ;
        RECT 1.485 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.170 ;
        RECT 0.340 -0.085 0.940 0.085 ;
        RECT 0.940 -0.085 1.305 0.170 ;
        RECT 1.305 -0.085 1.395 0.085 ;
        RECT 1.395 -0.085 1.485 0.490 ;
        RECT 1.485 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.320 ;
      RECT 0.220 0.410 0.300 1.090 ;
      RECT 0.300 1.005 0.390 1.090 ;
      RECT 0.125 0.250 0.430 0.320 ;
      RECT 0.390 1.005 0.495 1.245 ;
      RECT 0.430 0.175 0.550 0.320 ;
      RECT 0.300 0.410 0.640 0.490 ;
      RECT 0.640 0.175 0.730 0.490 ;
      RECT 0.525 0.870 0.905 0.940 ;
      RECT 0.905 0.655 0.985 0.940 ;
      RECT 0.495 1.005 1.070 1.080 ;
      RECT 1.070 0.825 1.150 1.080 ;
      RECT 0.585 1.145 1.150 1.225 ;
      RECT 0.985 0.655 1.215 0.735 ;
      RECT 1.215 0.385 1.305 1.225 ;
  END
END ACELEM1X1

MACRO ACELEM1X2
  CLASS CORE ;
  FOREIGN ACELEM1X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.595 0.845 0.805 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.420 0.130 1.015 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.935 0.595 1.150 0.805 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.175 1.665 1.150 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.105 0.130 1.485 ;
        RECT 0.130 1.315 0.795 1.485 ;
        RECT 0.795 1.240 0.940 1.485 ;
        RECT 0.940 1.315 1.395 1.485 ;
        RECT 1.395 0.895 1.485 1.485 ;
        RECT 1.485 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.170 ;
        RECT 0.340 -0.085 0.995 0.085 ;
        RECT 0.995 -0.085 1.125 0.205 ;
        RECT 1.125 -0.085 1.395 0.085 ;
        RECT 1.395 -0.085 1.485 0.230 ;
        RECT 1.485 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.115 0.330 ;
      RECT 0.220 0.420 0.290 1.225 ;
      RECT 0.115 0.260 0.445 0.330 ;
      RECT 0.290 1.060 0.510 1.225 ;
      RECT 0.445 0.175 0.550 0.330 ;
      RECT 0.290 0.420 0.640 0.505 ;
      RECT 0.640 0.175 0.745 0.505 ;
      RECT 0.600 1.060 1.125 1.150 ;
      RECT 0.745 0.295 1.130 0.505 ;
      RECT 0.500 0.895 1.215 0.970 ;
      RECT 1.215 0.895 1.220 1.170 ;
      RECT 1.220 0.175 1.305 1.170 ;
  END
END ACELEM1X2

MACRO ACELEM1X4
  CLASS CORE ;
  FOREIGN ACELEM1X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.735 0.960 0.815 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.130 0.665 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.455 1.150 0.665 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.490 0.500 1.580 0.760 ;
        RECT 1.580 0.230 1.670 1.090 ;
        RECT 1.670 0.230 1.675 0.645 ;
        RECT 1.675 0.555 1.765 0.645 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.050 1.485 ;
        RECT 0.050 1.055 0.140 1.485 ;
        RECT 0.140 1.315 0.790 1.485 ;
        RECT 0.790 1.240 0.930 1.485 ;
        RECT 0.930 1.315 1.400 1.485 ;
        RECT 1.400 0.860 1.490 1.485 ;
        RECT 1.490 1.315 1.765 1.485 ;
        RECT 1.765 0.735 1.855 1.485 ;
        RECT 1.855 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.210 0.085 ;
        RECT 0.210 -0.085 0.345 0.160 ;
        RECT 0.345 -0.085 1.005 0.085 ;
        RECT 1.005 -0.085 1.150 0.250 ;
        RECT 1.150 -0.085 1.400 0.085 ;
        RECT 1.400 -0.085 1.490 0.390 ;
        RECT 1.490 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.855 0.465 ;
        RECT 1.855 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.310 ;
      RECT 0.210 0.395 0.290 0.985 ;
      RECT 0.290 0.905 0.420 0.985 ;
      RECT 0.125 0.230 0.435 0.310 ;
      RECT 0.420 0.905 0.510 1.175 ;
      RECT 0.435 0.175 0.525 0.310 ;
      RECT 0.290 0.395 0.615 0.475 ;
      RECT 0.615 0.175 0.700 0.475 ;
      RECT 0.565 0.565 0.790 0.645 ;
      RECT 0.790 0.315 0.870 0.645 ;
      RECT 0.510 0.905 1.050 0.985 ;
      RECT 0.600 1.070 1.125 1.150 ;
      RECT 1.050 0.755 1.130 0.985 ;
      RECT 0.870 0.315 1.215 0.390 ;
      RECT 1.215 0.315 1.310 1.150 ;
  END
END ACELEM1X4

MACRO FILL1
  CLASS CORE SPACER ;
  FOREIGN FILL1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.190 BY 1.400 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.190 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.190 0.085 ;
    END
  END VSS
END FILL1

MACRO FILLTIE
  CLASS CORE WELLTAP ;
  FOREIGN FILLTIE 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.190 BY 1.400 ;
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.040 1.485 ;
        RECT 0.040 1.255 0.110 1.485 ;
        RECT 0.110 1.315 0.190 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.040 0.085 ;
        RECT 0.040 -0.085 0.110 0.145 ;
        RECT 0.110 -0.085 0.190 0.085 ;
    END
  END VSS
END FILLTIE

MACRO INCL1W1111OF4X1
  CLASS CORE ;
  FOREIGN INCL1W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.310 0.150 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.215 0.715 0.540 1.155 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.375 0.565 0.650 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.810 0.280 0.900 0.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.089600 ;
    PORT
      LAYER metal1 ;
        RECT 0.215 0.150 0.345 0.595 ;
        RECT 0.345 0.240 0.630 0.310 ;
        RECT 0.630 0.150 0.720 1.215 ;
        RECT 0.720 0.940 0.905 1.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.060 1.485 ;
        RECT 0.060 0.940 0.150 1.485 ;
        RECT 0.150 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.060 0.085 ;
        RECT 0.060 -0.085 0.150 0.240 ;
        RECT 0.150 -0.085 0.410 0.085 ;
        RECT 0.410 -0.085 0.560 0.175 ;
        RECT 0.560 -0.085 0.810 0.085 ;
        RECT 0.810 -0.085 0.905 0.215 ;
        RECT 0.905 -0.085 0.950 0.085 ;
    END
  END VSS
END INCL1W1111OF4X1

MACRO INCL1W111OF3X1
  CLASS CORE ;
  FOREIGN INCL1W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.385 0.145 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.375 0.730 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.800 0.755 1.060 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.125925 ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.150 0.335 1.225 ;
        RECT 0.335 1.150 0.820 1.225 ;
        RECT 0.820 0.150 0.905 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.055 1.485 ;
        RECT 0.055 0.940 0.180 1.485 ;
        RECT 0.180 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.055 0.085 ;
        RECT 0.055 -0.085 0.180 0.320 ;
        RECT 0.180 -0.085 0.440 0.085 ;
        RECT 0.440 -0.085 0.755 0.285 ;
        RECT 0.755 -0.085 0.950 0.085 ;
    END
  END VSS
END INCL1W111OF3X1

MACRO INCL1W11OF2X1
  CLASS CORE ;
  FOREIGN INCL1W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020250 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.320 0.510 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020250 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.320 0.160 0.875 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.049975 ;
    PORT
      LAYER metal1 ;
        RECT 0.250 0.180 0.340 1.225 ;
        RECT 0.340 0.940 0.525 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.070 1.485 ;
        RECT 0.070 0.940 0.160 1.485 ;
        RECT 0.160 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.070 0.085 ;
        RECT 0.070 -0.085 0.160 0.255 ;
        RECT 0.160 -0.085 0.420 0.085 ;
        RECT 0.420 -0.085 0.525 0.255 ;
        RECT 0.525 -0.085 0.570 0.085 ;
    END
  END VSS
END INCL1W11OF2X1

MACRO INCL1W11OF2X2
  CLASS CORE ;
  FOREIGN INCL1W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.040250 ;
    PORT
      LAYER metal1 ;
        RECT 0.425 0.365 0.515 0.740 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.040250 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.420 0.150 0.860 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.110200 ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.150 0.325 1.225 ;
        RECT 0.325 0.805 0.515 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.925 0.135 1.485 ;
        RECT 0.135 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.170 0.355 ;
        RECT 0.170 -0.085 0.390 0.085 ;
        RECT 0.390 -0.085 0.525 0.300 ;
        RECT 0.525 -0.085 0.570 0.085 ;
    END
  END VSS
END INCL1W11OF2X2

MACRO INCL1W1OF1X1
  CLASS CORE ;
  FOREIGN INCL1W1OF1X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.380 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.018000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.280 0.135 0.875 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.150 0.335 1.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.075 1.485 ;
        RECT 0.075 0.940 0.170 1.485 ;
        RECT 0.170 1.315 0.380 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.075 0.085 ;
        RECT 0.075 -0.085 0.175 0.215 ;
        RECT 0.175 -0.085 0.380 0.085 ;
    END
  END VSS
END INCL1W1OF1X1

MACRO INCL1W1OF1X2
  CLASS CORE ;
  FOREIGN INCL1W1OF1X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.380 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.036500 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.135 0.875 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.150 0.335 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.940 0.115 1.485 ;
        RECT 0.115 0.940 0.180 1.030 ;
        RECT 0.115 1.315 0.380 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.180 0.320 ;
        RECT 0.180 -0.085 0.380 0.085 ;
    END
  END VSS
END INCL1W1OF1X2

MACRO INCL1W1OF1X4
  CLASS CORE ;
  FOREIGN INCL1W1OF1X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.073000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.135 0.875 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.102200 ;
    PORT
      LAYER metal1 ;
        RECT 0.250 0.170 0.340 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.940 0.115 1.485 ;
        RECT 0.115 0.940 0.185 1.095 ;
        RECT 0.115 1.315 0.435 1.485 ;
        RECT 0.435 0.770 0.525 1.485 ;
        RECT 0.525 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.185 0.320 ;
        RECT 0.185 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.525 0.360 ;
        RECT 0.525 -0.085 0.570 0.085 ;
    END
  END VSS
END INCL1W1OF1X4

MACRO INCL2W11OF2X1
  CLASS CORE ;
  FOREIGN INCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.455 0.770 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.525 0.320 0.945 ;
        RECT 0.320 0.875 0.615 0.945 ;
        RECT 0.615 0.800 0.800 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.210 1.665 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.990 0.130 1.485 ;
        RECT 0.130 1.315 0.385 1.485 ;
        RECT 0.385 1.165 0.550 1.485 ;
        RECT 0.550 1.315 1.365 1.485 ;
        RECT 1.365 0.755 1.485 1.485 ;
        RECT 1.485 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.390 ;
        RECT 0.135 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.250 ;
        RECT 0.550 -0.085 1.350 0.085 ;
        RECT 1.350 -0.085 1.510 0.250 ;
        RECT 1.510 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200 0.315 0.615 0.390 ;
      RECT 0.200 1.010 0.615 1.100 ;
      RECT 0.615 0.175 0.685 0.390 ;
      RECT 0.615 1.010 0.700 1.225 ;
      RECT 0.775 0.310 0.865 0.390 ;
      RECT 0.865 0.310 0.945 1.090 ;
      RECT 0.945 0.310 0.965 0.525 ;
      RECT 0.700 1.155 1.010 1.225 ;
      RECT 0.685 0.175 1.030 0.245 ;
      RECT 1.030 0.175 1.120 0.385 ;
      RECT 1.185 0.210 1.275 0.385 ;
      RECT 1.035 0.590 1.275 0.935 ;
      RECT 1.010 1.000 1.300 1.225 ;
      RECT 0.965 0.450 1.345 0.525 ;
      RECT 1.275 0.315 1.420 0.385 ;
      RECT 1.275 0.590 1.420 0.680 ;
      RECT 1.420 0.315 1.510 0.680 ;
  END
END INCL2W11OF2X1

MACRO INCL2W11OF2X2
  CLASS CORE ;
  FOREIGN INCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.455 0.770 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.525 0.320 0.945 ;
        RECT 0.320 0.875 0.735 0.945 ;
        RECT 0.735 0.800 0.840 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.170 1.665 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.000 0.135 1.485 ;
        RECT 0.135 1.315 0.415 1.485 ;
        RECT 0.415 1.150 0.575 1.485 ;
        RECT 0.575 1.315 1.365 1.485 ;
        RECT 1.365 0.895 1.510 1.485 ;
        RECT 1.510 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.420 ;
        RECT 0.135 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.250 ;
        RECT 0.550 -0.085 1.375 0.085 ;
        RECT 1.375 -0.085 1.510 0.250 ;
        RECT 1.510 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200 0.315 0.615 0.390 ;
      RECT 0.200 1.010 0.640 1.085 ;
      RECT 0.615 0.175 0.685 0.390 ;
      RECT 0.640 1.010 0.710 1.225 ;
      RECT 0.815 0.315 0.905 0.405 ;
      RECT 0.905 0.315 0.980 1.085 ;
      RECT 0.685 0.175 1.045 0.250 ;
      RECT 0.710 1.150 1.045 1.225 ;
      RECT 1.045 0.175 1.155 0.420 ;
      RECT 1.045 0.945 1.300 1.225 ;
      RECT 1.220 0.150 1.310 0.420 ;
      RECT 0.980 0.495 1.375 0.605 ;
      RECT 1.310 0.315 1.440 0.420 ;
      RECT 1.045 0.695 1.440 0.830 ;
      RECT 1.440 0.315 1.510 0.830 ;
  END
END INCL2W11OF2X2

MACRO INCL2W11OF2X4
  CLASS CORE ;
  FOREIGN INCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042750 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.510 0.625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042750 ;
    PORT
      LAYER metal1 ;
        RECT 0.110 0.715 0.600 0.805 ;
        RECT 0.600 0.525 0.850 0.805 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.580 0.175 1.670 1.180 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.900 0.125 1.485 ;
        RECT 0.125 1.315 0.440 1.485 ;
        RECT 0.440 1.065 0.575 1.485 ;
        RECT 0.575 1.315 1.320 1.485 ;
        RECT 1.320 1.240 1.505 1.485 ;
        RECT 1.505 1.315 1.765 1.485 ;
        RECT 1.765 1.065 1.855 1.485 ;
        RECT 1.855 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.295 ;
        RECT 0.125 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.560 0.125 ;
        RECT 0.560 -0.085 1.395 0.085 ;
        RECT 1.395 -0.085 1.485 0.360 ;
        RECT 1.485 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.855 0.405 ;
        RECT 1.855 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 0.900 0.350 1.225 ;
      RECT 0.215 0.215 0.655 0.295 ;
      RECT 0.655 0.175 0.730 0.295 ;
      RECT 0.810 0.345 0.915 0.435 ;
      RECT 0.915 0.345 0.985 0.810 ;
      RECT 0.730 0.175 1.050 0.255 ;
      RECT 0.985 0.605 1.050 0.810 ;
      RECT 1.050 0.175 1.130 0.350 ;
      RECT 0.350 0.900 1.140 0.980 ;
      RECT 1.075 0.440 1.215 0.530 ;
      RECT 1.025 1.070 1.230 1.225 ;
      RECT 1.140 0.775 1.275 0.980 ;
      RECT 1.215 0.295 1.305 0.530 ;
      RECT 1.050 0.605 1.315 0.685 ;
      RECT 1.305 0.450 1.415 0.530 ;
      RECT 1.230 1.070 1.415 1.150 ;
      RECT 1.415 0.450 1.505 1.150 ;
  END
END INCL2W11OF2X4

MACRO INCL2W211OF3X1
  CLASS CORE ;
  FOREIGN INCL2W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024750 ;
    PORT
      LAYER metal1 ;
        RECT 1.390 0.245 1.475 0.455 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.095 0.595 0.580 0.810 ;
        RECT 0.580 0.720 0.710 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.310 0.455 0.800 0.530 ;
        RECT 0.800 0.455 0.890 0.735 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 1.915 0.220 1.955 0.480 ;
        RECT 1.955 0.220 2.045 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.970 0.135 1.485 ;
        RECT 0.135 1.315 0.405 1.485 ;
        RECT 0.405 1.070 0.540 1.485 ;
        RECT 0.540 1.315 1.705 1.485 ;
        RECT 1.705 1.210 1.860 1.485 ;
        RECT 1.860 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.310 ;
        RECT 0.135 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.540 0.195 ;
        RECT 0.540 -0.085 1.415 0.085 ;
        RECT 1.415 -0.085 1.550 0.160 ;
        RECT 1.550 -0.085 1.735 0.085 ;
        RECT 1.735 -0.085 1.825 0.455 ;
        RECT 1.825 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.195 0.315 0.365 ;
      RECT 0.225 0.900 0.315 1.225 ;
      RECT 0.315 0.285 0.630 0.365 ;
      RECT 0.315 0.900 0.630 0.980 ;
      RECT 0.630 0.175 0.710 0.365 ;
      RECT 0.630 0.900 0.710 1.225 ;
      RECT 0.800 0.310 0.955 0.390 ;
      RECT 0.955 0.310 1.035 0.820 ;
      RECT 0.710 0.175 1.100 0.245 ;
      RECT 1.100 0.175 1.180 0.310 ;
      RECT 0.710 1.135 1.200 1.225 ;
      RECT 1.035 0.400 1.245 0.480 ;
      RECT 0.800 0.910 1.320 1.045 ;
      RECT 1.245 0.175 1.325 0.480 ;
      RECT 1.035 0.740 1.415 0.820 ;
      RECT 1.125 0.570 1.565 0.650 ;
      RECT 1.410 1.040 1.615 1.225 ;
      RECT 1.565 0.400 1.645 0.650 ;
      RECT 1.415 0.740 1.690 0.945 ;
      RECT 1.645 0.560 1.780 0.650 ;
      RECT 1.615 1.040 1.780 1.120 ;
      RECT 1.780 0.560 1.865 1.120 ;
  END
END INCL2W211OF3X1

MACRO INCL2W211OF3X2
  CLASS CORE ;
  FOREIGN INCL2W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024750 ;
    PORT
      LAYER metal1 ;
        RECT 1.510 0.455 1.720 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.735 0.370 0.870 ;
        RECT 0.370 0.735 0.585 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.325 0.575 0.675 0.665 ;
        RECT 0.675 0.575 0.960 0.805 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.045 1.220 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.075 1.485 ;
        RECT 0.075 0.970 0.165 1.485 ;
        RECT 0.165 1.315 0.480 1.485 ;
        RECT 0.480 1.190 0.570 1.485 ;
        RECT 0.570 1.315 1.770 1.485 ;
        RECT 1.770 1.140 1.870 1.485 ;
        RECT 1.870 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.080 0.085 ;
        RECT 0.080 -0.085 0.170 0.315 ;
        RECT 0.170 -0.085 0.480 0.085 ;
        RECT 0.480 -0.085 0.570 0.315 ;
        RECT 0.570 -0.085 1.410 0.085 ;
        RECT 1.410 -0.085 1.515 0.210 ;
        RECT 1.515 -0.085 1.770 0.085 ;
        RECT 1.770 -0.085 1.870 0.210 ;
        RECT 1.870 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.260 0.260 0.355 0.485 ;
      RECT 0.255 1.020 0.390 1.225 ;
      RECT 0.355 0.405 0.660 0.485 ;
      RECT 0.390 1.020 0.660 1.100 ;
      RECT 0.660 0.175 0.740 0.485 ;
      RECT 0.660 1.020 0.740 1.225 ;
      RECT 0.830 0.330 0.970 0.485 ;
      RECT 0.970 0.405 1.025 0.485 ;
      RECT 0.740 0.175 1.050 0.255 ;
      RECT 1.025 0.405 1.095 0.805 ;
      RECT 1.050 0.175 1.130 0.315 ;
      RECT 0.740 1.145 1.165 1.225 ;
      RECT 1.095 0.720 1.185 0.805 ;
      RECT 1.095 0.405 1.205 0.485 ;
      RECT 1.205 0.175 1.285 0.485 ;
      RECT 1.185 0.720 1.320 0.925 ;
      RECT 1.160 0.550 1.350 0.630 ;
      RECT 0.830 1.000 1.410 1.080 ;
      RECT 1.350 0.300 1.430 0.630 ;
      RECT 1.410 0.925 1.490 1.080 ;
      RECT 1.580 0.970 1.680 1.150 ;
      RECT 1.320 0.755 1.705 0.835 ;
      RECT 1.430 0.300 1.795 0.380 ;
      RECT 1.680 0.970 1.795 1.050 ;
      RECT 1.795 0.300 1.875 1.050 ;
  END
END INCL2W211OF3X2

MACRO INCL2W211OF3X4
  CLASS CORE ;
  FOREIGN INCL2W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.575 1.395 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.100 0.735 0.370 0.825 ;
        RECT 0.370 0.735 0.635 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.345 0.455 0.845 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105125 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.050 1.125 ;
        RECT 2.050 0.560 2.140 0.665 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.125 1.485 ;
        RECT 0.125 1.315 0.430 1.485 ;
        RECT 0.430 1.190 0.520 1.485 ;
        RECT 0.520 1.315 1.775 1.485 ;
        RECT 1.775 1.050 1.870 1.485 ;
        RECT 1.870 1.315 2.140 1.485 ;
        RECT 2.140 0.910 2.230 1.485 ;
        RECT 2.230 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.195 ;
        RECT 0.135 -0.085 0.430 0.085 ;
        RECT 0.430 -0.085 0.520 0.195 ;
        RECT 0.520 -0.085 1.435 0.085 ;
        RECT 1.435 -0.085 1.655 0.225 ;
        RECT 1.655 -0.085 1.775 0.085 ;
        RECT 1.775 -0.085 1.870 0.495 ;
        RECT 1.870 -0.085 2.140 0.085 ;
        RECT 2.140 -0.085 2.230 0.470 ;
        RECT 2.230 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.175 0.340 0.365 ;
      RECT 0.205 1.020 0.340 1.225 ;
      RECT 0.340 0.285 0.610 0.365 ;
      RECT 0.340 1.020 0.610 1.100 ;
      RECT 0.610 0.175 0.700 0.365 ;
      RECT 0.610 1.020 0.700 1.225 ;
      RECT 0.790 0.310 0.915 0.390 ;
      RECT 0.915 0.310 0.995 0.935 ;
      RECT 0.700 0.175 1.085 0.245 ;
      RECT 0.700 1.145 1.130 1.225 ;
      RECT 1.085 0.175 1.165 0.315 ;
      RECT 0.995 0.405 1.255 0.485 ;
      RECT 0.790 1.000 1.285 1.080 ;
      RECT 1.255 0.175 1.345 0.485 ;
      RECT 0.995 0.865 1.375 0.935 ;
      RECT 1.085 0.730 1.515 0.800 ;
      RECT 1.375 0.865 1.515 1.225 ;
      RECT 1.515 0.400 1.605 0.800 ;
      RECT 1.580 0.985 1.605 1.185 ;
      RECT 1.605 0.585 1.685 1.185 ;
      RECT 1.685 0.585 1.875 0.860 ;
  END
END INCL2W211OF3X4

MACRO INCL3W111OF3X1
  CLASS CORE ;
  FOREIGN INCL3W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.655 0.595 1.595 0.665 ;
        RECT 1.595 0.360 1.740 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.730 1.720 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047750 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.445 1.530 0.530 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 1.870 0.225 1.960 0.395 ;
        RECT 1.960 0.225 2.045 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.215 1.485 ;
        RECT 0.215 0.875 0.305 1.485 ;
        RECT 0.305 1.315 1.705 1.485 ;
        RECT 1.705 1.010 1.840 1.485 ;
        RECT 1.840 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.315 0.085 ;
        RECT 0.315 -0.085 0.465 0.335 ;
        RECT 0.465 -0.085 1.595 0.085 ;
        RECT 1.595 -0.085 1.805 0.290 ;
        RECT 1.805 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.245 0.115 1.015 ;
      RECT 0.115 0.740 0.150 1.015 ;
      RECT 0.115 0.245 0.250 0.335 ;
      RECT 0.150 0.740 0.370 0.810 ;
      RECT 0.370 0.740 0.440 1.225 ;
      RECT 0.180 0.400 0.505 0.675 ;
      RECT 0.505 0.400 0.585 0.945 ;
      RECT 0.535 0.175 0.625 0.335 ;
      RECT 0.585 0.400 0.695 0.530 ;
      RECT 0.695 0.310 0.800 0.530 ;
      RECT 0.625 0.175 1.060 0.245 ;
      RECT 0.505 1.010 1.060 1.090 ;
      RECT 0.800 0.310 1.125 0.380 ;
      RECT 0.585 0.875 1.250 0.945 ;
      RECT 1.125 0.220 1.275 0.380 ;
      RECT 0.440 1.155 1.565 1.225 ;
      RECT 1.565 0.875 1.635 1.225 ;
      RECT 1.635 0.875 1.805 0.945 ;
      RECT 1.805 0.570 1.895 0.945 ;
  END
END INCL3W111OF3X1

MACRO INCL3W111OF3X2
  CLASS CORE ;
  FOREIGN INCL3W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.675 0.590 0.810 0.805 ;
        RECT 0.810 0.735 1.910 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.870 1.370 0.945 ;
        RECT 1.370 0.870 1.600 1.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.585 1.530 0.670 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.700 0.870 1.975 1.155 ;
        RECT 1.975 0.150 2.045 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 0.995 0.340 1.485 ;
        RECT 0.340 1.315 1.655 1.485 ;
        RECT 1.655 1.220 1.885 1.485 ;
        RECT 1.885 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.335 0.250 ;
        RECT 0.335 -0.085 1.655 0.085 ;
        RECT 1.655 -0.085 1.885 0.385 ;
        RECT 1.885 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.135 1.235 ;
      RECT 0.135 0.655 0.340 0.930 ;
      RECT 0.200 0.315 0.405 0.590 ;
      RECT 0.405 0.315 0.475 1.080 ;
      RECT 0.540 0.450 0.610 0.895 ;
      RECT 0.400 0.175 1.105 0.250 ;
      RECT 0.445 1.145 1.105 1.225 ;
      RECT 0.475 0.315 1.170 0.385 ;
      RECT 0.475 1.010 1.170 1.080 ;
      RECT 1.170 0.225 1.305 0.385 ;
      RECT 1.170 1.010 1.305 1.250 ;
      RECT 0.610 0.450 1.655 0.520 ;
      RECT 1.655 0.450 1.910 0.670 ;
  END
END INCL3W111OF3X2

MACRO INCL3W111OF3X4
  CLASS CORE ;
  FOREIGN INCL3W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.610 0.660 0.895 ;
        RECT 0.660 0.610 0.755 0.805 ;
        RECT 0.755 0.730 1.720 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.870 1.530 0.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.585 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105125 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.050 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.265 1.485 ;
        RECT 0.265 0.955 0.355 1.485 ;
        RECT 0.355 1.315 1.565 1.485 ;
        RECT 1.565 1.185 1.720 1.485 ;
        RECT 1.720 1.315 2.145 1.485 ;
        RECT 2.145 0.705 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.215 ;
        RECT 0.340 -0.085 1.565 0.085 ;
        RECT 1.565 -0.085 1.850 0.215 ;
        RECT 1.850 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.400 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.115 1.230 ;
      RECT 0.115 0.655 0.135 1.230 ;
      RECT 0.180 0.310 0.260 0.585 ;
      RECT 0.135 0.655 0.340 0.735 ;
      RECT 0.340 0.450 0.430 0.735 ;
      RECT 0.445 0.985 0.550 1.225 ;
      RECT 0.430 0.175 0.985 0.245 ;
      RECT 0.550 1.155 1.035 1.225 ;
      RECT 0.260 0.310 1.075 0.385 ;
      RECT 1.075 0.210 1.250 0.385 ;
      RECT 0.430 0.450 1.625 0.520 ;
      RECT 1.625 0.450 1.750 0.615 ;
      RECT 1.250 0.305 1.815 0.385 ;
      RECT 0.640 1.015 1.815 1.090 ;
      RECT 1.815 0.305 1.895 1.090 ;
  END
END INCL3W111OF3X4

MACRO INCL3W211OF3X1
  CLASS CORE ;
  FOREIGN INCL3W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.970 0.595 1.465 0.680 ;
        RECT 1.465 0.595 1.650 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.870 0.560 0.960 ;
        RECT 0.560 0.550 0.770 0.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.455 0.390 0.805 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.245 2.235 1.015 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.410 1.485 ;
        RECT 0.410 1.225 0.635 1.485 ;
        RECT 0.635 1.315 1.545 1.485 ;
        RECT 1.545 1.095 1.680 1.485 ;
        RECT 1.680 1.315 1.915 1.485 ;
        RECT 1.915 0.710 2.055 1.485 ;
        RECT 2.055 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.065 0.085 ;
        RECT 0.065 -0.085 0.155 0.280 ;
        RECT 0.155 -0.085 0.410 0.085 ;
        RECT 0.410 -0.085 0.565 0.245 ;
        RECT 0.565 -0.085 0.790 0.085 ;
        RECT 0.790 -0.085 0.975 0.110 ;
        RECT 0.975 -0.085 1.915 0.085 ;
        RECT 1.915 -0.085 2.060 0.305 ;
        RECT 2.060 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235 0.215 0.325 0.390 ;
      RECT 0.045 1.045 0.700 1.135 ;
      RECT 0.700 1.045 0.770 1.225 ;
      RECT 0.835 0.455 0.905 0.850 ;
      RECT 0.905 0.780 1.015 0.850 ;
      RECT 0.325 0.310 1.200 0.390 ;
      RECT 1.015 0.780 1.200 1.070 ;
      RECT 0.905 0.455 1.350 0.530 ;
      RECT 1.265 0.745 1.400 1.010 ;
      RECT 0.770 1.135 1.480 1.225 ;
      RECT 1.350 0.310 1.485 0.530 ;
      RECT 0.630 0.175 1.550 0.245 ;
      RECT 1.550 0.175 1.655 0.330 ;
      RECT 1.485 0.395 1.695 0.530 ;
      RECT 1.400 0.940 1.760 1.010 ;
      RECT 1.760 0.245 1.845 1.010 ;
      RECT 1.845 0.245 1.850 0.645 ;
      RECT 1.850 0.370 2.060 0.645 ;
  END
END INCL3W211OF3X1

MACRO INCL3W211OF3X2
  CLASS CORE ;
  FOREIGN INCL3W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044500 ;
    PORT
      LAYER metal1 ;
        RECT 1.025 0.735 1.720 0.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.870 0.600 0.960 ;
        RECT 0.600 0.465 0.800 0.960 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.465 0.510 0.780 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078650 ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.150 2.235 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.425 1.485 ;
        RECT 0.425 1.170 0.590 1.485 ;
        RECT 0.590 1.315 1.580 1.485 ;
        RECT 1.580 1.070 1.720 1.485 ;
        RECT 1.720 1.315 1.945 1.485 ;
        RECT 1.945 0.870 2.040 1.485 ;
        RECT 2.040 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.055 0.085 ;
        RECT 0.055 -0.085 0.145 0.360 ;
        RECT 0.145 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.555 0.245 ;
        RECT 0.555 -0.085 0.790 0.085 ;
        RECT 0.790 -0.085 0.975 0.110 ;
        RECT 0.975 -0.085 1.910 0.085 ;
        RECT 1.910 -0.085 2.040 0.210 ;
        RECT 2.040 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 1.035 0.265 1.245 ;
      RECT 0.245 0.215 0.335 0.400 ;
      RECT 0.265 1.035 0.660 1.105 ;
      RECT 0.660 1.035 0.730 1.225 ;
      RECT 0.890 0.580 0.960 1.070 ;
      RECT 0.960 0.885 1.185 1.070 ;
      RECT 0.335 0.310 1.330 0.400 ;
      RECT 0.960 0.580 1.420 0.670 ;
      RECT 1.420 0.310 1.515 0.670 ;
      RECT 0.730 1.135 1.515 1.225 ;
      RECT 0.620 0.175 1.590 0.245 ;
      RECT 1.590 0.175 1.690 0.375 ;
      RECT 1.250 0.885 1.785 0.975 ;
      RECT 1.755 0.150 1.845 0.360 ;
      RECT 1.785 0.735 1.880 0.975 ;
      RECT 1.515 0.465 1.910 0.670 ;
      RECT 1.845 0.280 1.990 0.360 ;
      RECT 1.880 0.735 1.990 0.805 ;
      RECT 1.990 0.280 2.080 0.805 ;
  END
END INCL3W211OF3X2

MACRO INCL3W211OF3X4
  CLASS CORE ;
  FOREIGN INCL3W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.980 0.525 1.135 0.945 ;
        RECT 1.135 0.855 1.565 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.715 0.350 0.945 ;
        RECT 0.350 0.855 0.865 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.320 0.525 0.440 0.615 ;
        RECT 0.440 0.525 0.890 0.765 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.124100 ;
    PORT
      LAYER metal1 ;
        RECT 2.275 0.185 2.410 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.425 1.485 ;
        RECT 0.425 1.240 0.585 1.485 ;
        RECT 0.585 1.315 1.620 1.485 ;
        RECT 1.620 1.205 1.725 1.485 ;
        RECT 1.725 1.315 2.050 1.485 ;
        RECT 2.050 1.025 2.185 1.485 ;
        RECT 2.185 1.315 2.500 1.485 ;
        RECT 2.500 0.870 2.580 1.485 ;
        RECT 2.580 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.170 0.305 ;
        RECT 0.170 -0.085 0.440 0.085 ;
        RECT 0.440 -0.085 0.540 0.265 ;
        RECT 0.540 -0.085 0.855 0.085 ;
        RECT 0.855 -0.085 1.010 0.110 ;
        RECT 1.010 -0.085 2.050 0.085 ;
        RECT 2.050 -0.085 2.185 0.415 ;
        RECT 2.185 -0.085 2.500 0.085 ;
        RECT 2.500 -0.085 2.580 0.420 ;
        RECT 2.580 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.260 0.185 0.350 0.435 ;
      RECT 0.060 1.035 0.675 1.170 ;
      RECT 0.675 1.035 0.745 1.225 ;
      RECT 0.350 0.355 1.195 0.435 ;
      RECT 1.260 0.355 1.330 0.765 ;
      RECT 0.745 1.145 1.530 1.225 ;
      RECT 1.330 0.355 1.535 0.435 ;
      RECT 0.630 0.185 1.645 0.265 ;
      RECT 1.330 0.685 1.655 0.765 ;
      RECT 1.050 1.010 1.655 1.080 ;
      RECT 1.645 0.185 1.735 0.420 ;
      RECT 1.655 0.685 1.735 1.080 ;
      RECT 1.395 0.525 1.825 0.605 ;
      RECT 1.825 0.385 1.960 0.605 ;
      RECT 1.825 0.855 1.960 1.085 ;
      RECT 1.735 0.685 2.015 0.765 ;
      RECT 1.960 0.505 2.105 0.605 ;
      RECT 1.960 0.855 2.105 0.935 ;
      RECT 2.105 0.505 2.185 0.935 ;
  END
END INCL3W211OF3X4

MACRO INCL4W1111OF4X1
  CLASS CORE ;
  FOREIGN INCL4W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.550 0.425 0.850 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.450 0.480 0.805 ;
        RECT 0.480 0.730 1.040 0.805 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.395 1.105 0.665 ;
        RECT 0.180 0.870 1.105 0.960 ;
        RECT 1.105 0.395 1.195 0.960 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.395 0.500 1.775 0.775 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.235 2.240 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.230 1.485 ;
        RECT 0.230 1.180 0.385 1.485 ;
        RECT 0.385 1.315 0.590 1.485 ;
        RECT 0.590 1.180 0.755 1.485 ;
        RECT 0.755 1.315 1.760 1.485 ;
        RECT 1.760 0.975 1.895 1.485 ;
        RECT 1.895 1.315 2.335 1.485 ;
        RECT 2.335 0.680 2.425 1.485 ;
        RECT 2.425 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.365 0.225 ;
        RECT 0.365 -0.085 0.590 0.085 ;
        RECT 0.590 -0.085 0.745 0.225 ;
        RECT 0.745 -0.085 1.795 0.085 ;
        RECT 1.795 -0.085 1.930 0.275 ;
        RECT 1.930 -0.085 2.335 0.085 ;
        RECT 2.335 -0.085 2.425 0.495 ;
        RECT 2.425 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.165 0.135 0.360 ;
      RECT 0.135 0.290 0.435 0.360 ;
      RECT 0.435 0.165 0.525 0.360 ;
      RECT 0.525 0.290 0.810 0.360 ;
      RECT 0.045 1.025 0.825 1.115 ;
      RECT 0.810 0.175 0.880 0.360 ;
      RECT 0.825 1.025 0.895 1.225 ;
      RECT 1.260 0.310 1.330 1.080 ;
      RECT 1.330 0.975 1.505 1.080 ;
      RECT 1.330 0.310 1.510 0.410 ;
      RECT 0.880 0.175 1.570 0.245 ;
      RECT 0.895 1.145 1.570 1.225 ;
      RECT 1.570 0.975 1.695 1.225 ;
      RECT 1.570 0.175 1.730 0.275 ;
      RECT 1.510 0.340 1.840 0.410 ;
      RECT 1.840 0.340 1.930 0.695 ;
      RECT 1.490 0.840 1.995 0.910 ;
      RECT 1.995 0.235 2.085 1.250 ;
  END
END INCL4W1111OF4X1

MACRO INCL4W1111OF4X2
  CLASS CORE ;
  FOREIGN INCL4W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.350 0.595 0.650 0.810 ;
        RECT 0.650 0.595 0.835 0.685 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.325 0.435 0.900 0.525 ;
        RECT 0.900 0.435 1.025 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.260 0.965 ;
        RECT 0.260 0.875 1.090 0.965 ;
        RECT 1.090 0.535 1.180 0.965 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 1.380 0.535 1.465 0.875 ;
        RECT 1.465 0.805 1.580 0.875 ;
        RECT 1.580 0.805 1.715 1.015 ;
        RECT 1.715 0.805 1.815 0.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.805 2.335 1.105 ;
        RECT 2.335 0.195 2.425 1.105 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.225 0.355 1.485 ;
        RECT 0.355 1.315 0.580 1.485 ;
        RECT 0.580 1.225 0.780 1.485 ;
        RECT 0.780 1.315 1.780 1.485 ;
        RECT 1.780 0.940 1.915 1.485 ;
        RECT 1.915 1.315 2.150 1.485 ;
        RECT 2.150 1.170 2.265 1.485 ;
        RECT 2.265 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.170 ;
        RECT 0.355 -0.085 0.580 0.085 ;
        RECT 0.580 -0.085 0.780 0.170 ;
        RECT 0.780 -0.085 1.780 0.085 ;
        RECT 1.780 -0.085 1.915 0.335 ;
        RECT 1.915 -0.085 2.165 0.085 ;
        RECT 2.165 -0.085 2.265 0.400 ;
        RECT 2.265 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.140 0.305 ;
      RECT 0.045 1.080 0.140 1.250 ;
      RECT 0.140 0.235 0.425 0.305 ;
      RECT 0.425 0.150 0.515 0.305 ;
      RECT 1.245 0.370 1.315 1.015 ;
      RECT 1.315 0.370 1.515 0.470 ;
      RECT 1.315 0.940 1.515 1.015 ;
      RECT 0.515 0.235 1.575 0.305 ;
      RECT 1.530 0.535 1.670 0.740 ;
      RECT 1.575 0.235 1.715 0.335 ;
      RECT 0.140 1.080 1.715 1.160 ;
      RECT 1.515 0.400 1.810 0.470 ;
      RECT 1.810 0.400 1.915 0.595 ;
      RECT 1.670 0.660 1.995 0.740 ;
      RECT 1.995 0.300 2.085 1.180 ;
      RECT 2.085 0.300 2.100 0.730 ;
      RECT 2.100 0.465 2.265 0.730 ;
  END
END INCL4W1111OF4X2

MACRO INCL4W1111OF4X4
  CLASS CORE ;
  FOREIGN INCL4W1111OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.435 0.770 0.640 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.730 0.915 0.810 ;
        RECT 0.915 0.435 1.010 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.140 0.730 0.275 0.950 ;
        RECT 0.275 0.875 1.100 0.950 ;
        RECT 1.100 0.645 1.190 0.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.390 0.590 1.510 0.725 ;
        RECT 1.510 0.590 1.720 0.805 ;
        RECT 1.720 0.590 1.910 0.665 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 2.340 0.220 2.430 1.085 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.240 0.375 1.485 ;
        RECT 0.375 1.315 0.590 1.485 ;
        RECT 0.590 1.240 0.815 1.485 ;
        RECT 0.815 1.315 1.810 1.485 ;
        RECT 1.810 1.035 1.900 1.485 ;
        RECT 1.900 1.315 2.160 1.485 ;
        RECT 2.160 0.730 2.250 1.485 ;
        RECT 2.250 1.315 2.525 1.485 ;
        RECT 2.525 0.730 2.615 1.485 ;
        RECT 2.615 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.175 ;
        RECT 0.340 -0.085 0.590 0.085 ;
        RECT 0.590 -0.085 0.785 0.175 ;
        RECT 0.785 -0.085 1.790 0.085 ;
        RECT 1.790 -0.085 1.880 0.350 ;
        RECT 1.880 -0.085 2.160 0.085 ;
        RECT 2.160 -0.085 2.250 0.405 ;
        RECT 2.250 -0.085 2.525 0.085 ;
        RECT 2.525 -0.085 2.615 0.440 ;
        RECT 2.615 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.345 ;
      RECT 0.125 0.265 0.430 0.345 ;
      RECT 0.430 0.175 0.510 0.345 ;
      RECT 0.510 0.265 0.875 0.345 ;
      RECT 0.875 0.175 1.010 0.345 ;
      RECT 1.255 0.310 1.325 0.950 ;
      RECT 1.325 0.310 1.520 0.390 ;
      RECT 1.010 0.175 1.610 0.245 ;
      RECT 1.610 0.175 1.700 0.350 ;
      RECT 0.045 1.040 1.720 1.175 ;
      RECT 1.325 0.870 1.825 0.950 ;
      RECT 1.825 0.730 1.915 0.950 ;
      RECT 1.510 0.455 1.980 0.525 ;
      RECT 1.980 0.265 2.000 0.525 ;
      RECT 2.000 0.265 2.070 1.175 ;
      RECT 2.070 0.495 2.080 1.175 ;
      RECT 2.080 0.495 2.250 0.640 ;
  END
END INCL4W1111OF4X4

MACRO INCLP1W1111OF4X1
  CLASS CORE ;
  FOREIGN INCLP1W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024250 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.525 0.350 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024250 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.245 0.510 0.455 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024250 ;
    PORT
      LAYER metal1 ;
        RECT 0.575 0.245 0.710 0.595 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024250 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.665 0.770 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.095850 ;
    PORT
      LAYER metal1 ;
        RECT 0.800 0.220 0.835 0.455 ;
        RECT 0.235 1.035 0.835 1.130 ;
        RECT 0.835 0.220 0.905 1.130 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.055 1.485 ;
        RECT 0.055 1.060 0.145 1.485 ;
        RECT 0.145 1.315 0.405 1.485 ;
        RECT 0.405 1.220 0.555 1.485 ;
        RECT 0.555 1.315 0.775 1.485 ;
        RECT 0.775 1.205 0.905 1.485 ;
        RECT 0.905 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.200 0.160 ;
        RECT 0.200 -0.085 0.950 0.085 ;
    END
  END VSS
END INCLP1W1111OF4X1

MACRO INCLP1W111OF3X1
  CLASS CORE ;
  FOREIGN INCLP1W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.245 0.535 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.320 0.855 0.600 0.945 ;
        RECT 0.600 0.665 0.890 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.385 0.905 0.600 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.084925 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.165 0.255 1.245 ;
        RECT 0.255 1.010 0.350 1.245 ;
        RECT 0.350 1.010 0.905 1.085 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.975 0.115 1.485 ;
        RECT 0.115 1.315 0.420 1.485 ;
        RECT 0.420 1.150 0.695 1.485 ;
        RECT 0.695 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.690 0.085 ;
        RECT 0.690 -0.085 0.860 0.320 ;
        RECT 0.860 -0.085 0.950 0.085 ;
    END
  END VSS
END INCLP1W111OF3X1

MACRO INCLP1W11OF2X1
  CLASS CORE ;
  FOREIGN INCLP1W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.245 0.355 0.745 ;
        RECT 0.355 0.335 0.445 0.630 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.330 0.135 0.875 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.158475 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.155 0.510 0.270 ;
        RECT 0.235 0.875 0.510 1.175 ;
        RECT 0.510 0.155 0.580 1.175 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.080 1.485 ;
        RECT 0.080 0.940 0.170 1.485 ;
        RECT 0.170 1.315 0.645 1.485 ;
        RECT 0.645 0.615 0.715 1.485 ;
        RECT 0.715 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.080 0.085 ;
        RECT 0.080 -0.085 0.170 0.265 ;
        RECT 0.170 -0.085 0.760 0.085 ;
    END
  END VSS
END INCLP1W11OF2X1

MACRO INCLP1W11OF2X2
  CLASS CORE ;
  FOREIGN INCLP1W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.038750 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.520 0.510 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.038750 ;
    PORT
      LAYER metal1 ;
        RECT 0.050 0.385 0.140 0.745 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.097700 ;
    PORT
      LAYER metal1 ;
        RECT 0.245 0.155 0.335 1.195 ;
        RECT 0.335 0.155 0.525 0.455 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.075 1.485 ;
        RECT 0.075 0.810 0.165 1.485 ;
        RECT 0.165 1.315 0.435 1.485 ;
        RECT 0.435 0.940 0.525 1.485 ;
        RECT 0.525 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.180 0.320 ;
        RECT 0.180 -0.085 0.570 0.085 ;
    END
  END VSS
END INCLP1W11OF2X2

MACRO INCLP2W11OF2X1
  CLASS CORE ;
  FOREIGN INCLP2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.455 0.770 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.525 0.320 0.945 ;
        RECT 0.320 0.875 0.615 0.945 ;
        RECT 0.615 0.800 0.800 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.210 1.665 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.990 0.130 1.485 ;
        RECT 0.130 1.315 0.385 1.485 ;
        RECT 0.385 1.165 0.550 1.485 ;
        RECT 0.550 1.315 1.365 1.485 ;
        RECT 1.365 0.755 1.485 1.485 ;
        RECT 1.485 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.390 ;
        RECT 0.135 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.250 ;
        RECT 0.550 -0.085 1.350 0.085 ;
        RECT 1.350 -0.085 1.510 0.250 ;
        RECT 1.510 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200 0.315 0.615 0.390 ;
      RECT 0.200 1.010 0.615 1.100 ;
      RECT 0.615 0.175 0.685 0.390 ;
      RECT 0.615 1.010 0.700 1.225 ;
      RECT 0.775 0.310 0.865 0.390 ;
      RECT 0.865 0.310 0.945 1.090 ;
      RECT 0.945 0.310 0.965 0.525 ;
      RECT 0.700 1.155 1.010 1.225 ;
      RECT 0.685 0.175 1.030 0.245 ;
      RECT 1.030 0.175 1.120 0.385 ;
      RECT 1.185 0.210 1.275 0.385 ;
      RECT 1.035 0.590 1.275 0.935 ;
      RECT 1.010 1.000 1.300 1.225 ;
      RECT 0.965 0.450 1.345 0.525 ;
      RECT 1.275 0.315 1.420 0.385 ;
      RECT 1.275 0.590 1.420 0.680 ;
      RECT 1.420 0.315 1.510 0.680 ;
  END
END INCLP2W11OF2X1

MACRO INCLP2W11OF2X2
  CLASS CORE ;
  FOREIGN INCLP2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.385 0.455 0.770 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.525 0.320 0.945 ;
        RECT 0.320 0.875 0.735 0.945 ;
        RECT 0.735 0.800 0.840 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 1.575 0.170 1.665 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.000 0.135 1.485 ;
        RECT 0.135 1.315 0.415 1.485 ;
        RECT 0.415 1.150 0.575 1.485 ;
        RECT 0.575 1.315 1.365 1.485 ;
        RECT 1.365 0.895 1.510 1.485 ;
        RECT 1.510 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.420 ;
        RECT 0.135 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.250 ;
        RECT 0.550 -0.085 1.375 0.085 ;
        RECT 1.375 -0.085 1.510 0.250 ;
        RECT 1.510 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200 0.315 0.615 0.390 ;
      RECT 0.200 1.010 0.640 1.085 ;
      RECT 0.615 0.175 0.685 0.390 ;
      RECT 0.640 1.010 0.710 1.225 ;
      RECT 0.815 0.315 0.905 0.405 ;
      RECT 0.905 0.315 0.980 1.085 ;
      RECT 0.685 0.175 1.045 0.250 ;
      RECT 0.710 1.150 1.045 1.225 ;
      RECT 1.045 0.175 1.155 0.420 ;
      RECT 1.045 0.945 1.300 1.225 ;
      RECT 1.220 0.150 1.310 0.420 ;
      RECT 0.980 0.495 1.375 0.605 ;
      RECT 1.310 0.315 1.440 0.420 ;
      RECT 1.045 0.695 1.440 0.830 ;
      RECT 1.440 0.315 1.510 0.830 ;
  END
END INCLP2W11OF2X2

MACRO INCLP2W11OF2X4
  CLASS CORE ;
  FOREIGN INCLP2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.510 0.625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.110 0.715 0.600 0.805 ;
        RECT 0.600 0.525 0.850 0.805 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.580 0.175 1.670 1.180 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.895 0.125 1.485 ;
        RECT 0.125 1.315 0.440 1.485 ;
        RECT 0.440 1.065 0.575 1.485 ;
        RECT 0.575 1.315 1.320 1.485 ;
        RECT 1.320 1.235 1.500 1.485 ;
        RECT 1.500 1.315 1.765 1.485 ;
        RECT 1.765 1.065 1.855 1.485 ;
        RECT 1.855 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.295 ;
        RECT 0.125 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.575 0.125 ;
        RECT 0.575 -0.085 1.395 0.085 ;
        RECT 1.395 -0.085 1.495 0.360 ;
        RECT 1.495 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.855 0.405 ;
        RECT 1.855 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 0.895 0.350 1.225 ;
      RECT 0.215 0.215 0.655 0.295 ;
      RECT 0.655 0.175 0.730 0.295 ;
      RECT 0.810 0.345 0.915 0.435 ;
      RECT 0.915 0.345 0.985 0.805 ;
      RECT 0.730 0.175 1.050 0.255 ;
      RECT 0.985 0.600 1.050 0.805 ;
      RECT 1.050 0.175 1.130 0.350 ;
      RECT 0.350 0.895 1.140 0.975 ;
      RECT 1.075 0.440 1.215 0.530 ;
      RECT 1.025 1.065 1.230 1.225 ;
      RECT 1.140 0.770 1.275 0.975 ;
      RECT 1.215 0.295 1.305 0.530 ;
      RECT 1.050 0.600 1.325 0.680 ;
      RECT 1.305 0.450 1.415 0.530 ;
      RECT 1.230 1.065 1.415 1.145 ;
      RECT 1.415 0.450 1.505 1.145 ;
  END
END INCLP2W11OF2X4

MACRO INCLP2W211OF3X1
  CLASS CORE ;
  FOREIGN INCLP2W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 1.010 0.525 1.300 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.150 0.685 0.665 0.890 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.510 0.595 ;
        RECT 0.510 0.515 0.815 0.595 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.041800 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.385 2.235 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.980 0.125 1.485 ;
        RECT 0.125 1.315 0.415 1.485 ;
        RECT 0.415 1.150 0.560 1.485 ;
        RECT 0.560 1.315 1.520 1.485 ;
        RECT 1.520 1.290 1.700 1.485 ;
        RECT 1.700 1.315 1.960 1.485 ;
        RECT 1.960 1.090 2.050 1.485 ;
        RECT 2.050 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.295 ;
        RECT 0.125 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.560 0.125 ;
        RECT 0.560 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.050 0.430 ;
        RECT 2.050 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.205 0.215 0.650 0.295 ;
      RECT 0.205 0.980 0.650 1.060 ;
      RECT 0.650 0.175 0.730 0.295 ;
      RECT 0.650 0.980 0.730 1.225 ;
      RECT 0.820 0.330 0.965 0.425 ;
      RECT 0.730 0.175 1.160 0.255 ;
      RECT 0.730 1.135 1.160 1.225 ;
      RECT 0.965 0.345 1.225 0.425 ;
      RECT 1.225 0.215 1.305 0.425 ;
      RECT 0.820 0.965 1.390 1.045 ;
      RECT 1.390 0.385 1.480 1.045 ;
      RECT 1.480 0.690 1.490 1.045 ;
      RECT 1.305 0.215 1.570 0.295 ;
      RECT 1.570 0.215 1.660 0.520 ;
      RECT 1.235 1.120 1.750 1.200 ;
      RECT 1.750 0.385 1.870 0.600 ;
      RECT 1.750 0.920 1.870 1.200 ;
      RECT 1.490 0.690 1.895 0.785 ;
      RECT 1.870 0.520 1.985 0.600 ;
      RECT 1.870 0.920 1.985 1.000 ;
      RECT 1.985 0.520 2.065 1.000 ;
  END
END INCLP2W211OF3X1

MACRO INCLP2W211OF3X2
  CLASS CORE ;
  FOREIGN INCLP2W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022500 ;
    PORT
      LAYER metal1 ;
        RECT 1.200 0.595 1.575 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.130 0.735 0.585 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.315 0.585 0.690 0.665 ;
        RECT 0.690 0.585 0.960 0.805 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 2.005 0.800 2.145 0.945 ;
        RECT 2.145 0.800 2.150 1.170 ;
        RECT 2.150 0.175 2.235 1.170 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.065 0.125 1.485 ;
        RECT 0.125 1.315 0.410 1.485 ;
        RECT 0.410 1.225 0.545 1.485 ;
        RECT 0.545 1.315 1.535 1.485 ;
        RECT 1.535 1.260 1.675 1.485 ;
        RECT 1.675 1.315 1.800 1.485 ;
        RECT 1.800 1.240 2.060 1.485 ;
        RECT 2.060 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.055 0.085 ;
        RECT 0.055 -0.085 0.145 0.465 ;
        RECT 0.145 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.515 0.325 ;
        RECT 0.515 -0.085 1.800 0.085 ;
        RECT 1.800 -0.085 2.060 0.175 ;
        RECT 2.060 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.235 0.190 0.325 0.495 ;
      RECT 0.325 0.415 0.635 0.495 ;
      RECT 0.215 1.045 0.635 1.135 ;
      RECT 0.635 0.175 0.715 0.495 ;
      RECT 0.635 1.045 0.715 1.225 ;
      RECT 0.805 0.345 0.945 0.495 ;
      RECT 0.805 0.965 0.960 1.060 ;
      RECT 0.715 0.175 1.035 0.255 ;
      RECT 1.035 0.175 1.120 0.325 ;
      RECT 0.715 1.145 1.155 1.225 ;
      RECT 0.945 0.415 1.195 0.495 ;
      RECT 1.195 0.175 1.275 0.495 ;
      RECT 1.245 1.100 1.380 1.225 ;
      RECT 1.365 0.345 1.445 0.515 ;
      RECT 1.275 0.175 1.535 0.255 ;
      RECT 1.535 0.175 1.625 0.345 ;
      RECT 1.445 0.435 1.665 0.515 ;
      RECT 0.960 0.965 1.665 1.035 ;
      RECT 1.665 0.435 1.745 1.035 ;
      RECT 1.715 0.265 1.835 0.345 ;
      RECT 1.380 1.100 1.835 1.170 ;
      RECT 1.835 0.265 1.915 1.170 ;
      RECT 1.915 0.435 2.060 0.710 ;
  END
END INCLP2W211OF3X2

MACRO INCLP2W211OF3X4
  CLASS CORE ;
  FOREIGN INCLP2W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022250 ;
    PORT
      LAYER metal1 ;
        RECT 1.065 0.595 1.340 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.665 0.215 0.945 ;
        RECT 0.215 0.855 0.630 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.305 0.545 0.710 0.665 ;
        RECT 0.710 0.545 0.960 0.805 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105850 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.050 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.030 0.125 1.485 ;
        RECT 0.125 1.315 0.440 1.485 ;
        RECT 0.440 1.170 0.530 1.485 ;
        RECT 0.530 1.315 1.185 1.485 ;
        RECT 1.185 1.290 1.375 1.485 ;
        RECT 1.375 1.315 1.780 1.485 ;
        RECT 1.780 1.020 1.870 1.485 ;
        RECT 1.870 1.315 2.145 1.485 ;
        RECT 2.145 0.850 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.425 ;
        RECT 0.125 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.530 0.285 ;
        RECT 0.530 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.870 0.360 ;
        RECT 1.870 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.395 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.200 0.185 0.335 0.455 ;
      RECT 0.215 1.010 0.350 1.225 ;
      RECT 0.335 0.375 0.620 0.455 ;
      RECT 0.350 1.010 0.620 1.090 ;
      RECT 0.620 0.175 0.700 0.455 ;
      RECT 0.620 1.010 0.700 1.225 ;
      RECT 0.790 0.895 0.925 1.085 ;
      RECT 0.700 1.150 1.000 1.225 ;
      RECT 1.000 1.065 1.080 1.225 ;
      RECT 0.700 0.175 1.120 0.250 ;
      RECT 1.150 0.460 1.405 0.530 ;
      RECT 0.925 0.895 1.405 0.975 ;
      RECT 0.790 0.315 1.480 0.395 ;
      RECT 1.405 0.460 1.485 0.975 ;
      RECT 1.485 0.625 1.560 0.975 ;
      RECT 1.155 1.065 1.625 1.200 ;
      RECT 1.570 0.315 1.660 0.530 ;
      RECT 1.560 0.625 1.700 0.760 ;
      RECT 1.625 0.850 1.705 1.200 ;
      RECT 1.660 0.450 1.790 0.530 ;
      RECT 1.705 0.850 1.790 0.930 ;
      RECT 1.790 0.450 1.870 0.930 ;
  END
END INCLP2W211OF3X4

MACRO INCLP3W111OF3X1
  CLASS CORE ;
  FOREIGN INCLP3W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.655 0.595 1.595 0.665 ;
        RECT 1.595 0.360 1.740 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.730 1.720 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047750 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.445 1.530 0.530 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 1.870 0.225 1.960 0.395 ;
        RECT 1.960 0.225 2.045 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.215 1.485 ;
        RECT 0.215 0.875 0.305 1.485 ;
        RECT 0.305 1.315 1.705 1.485 ;
        RECT 1.705 1.010 1.840 1.485 ;
        RECT 1.840 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.315 0.085 ;
        RECT 0.315 -0.085 0.465 0.335 ;
        RECT 0.465 -0.085 1.595 0.085 ;
        RECT 1.595 -0.085 1.805 0.290 ;
        RECT 1.805 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.245 0.115 1.015 ;
      RECT 0.115 0.740 0.150 1.015 ;
      RECT 0.115 0.245 0.250 0.335 ;
      RECT 0.150 0.740 0.370 0.810 ;
      RECT 0.370 0.740 0.440 1.225 ;
      RECT 0.180 0.400 0.505 0.675 ;
      RECT 0.505 0.400 0.585 0.945 ;
      RECT 0.535 0.175 0.625 0.335 ;
      RECT 0.585 0.400 0.695 0.530 ;
      RECT 0.695 0.310 0.800 0.530 ;
      RECT 0.625 0.175 1.060 0.245 ;
      RECT 0.505 1.010 1.060 1.090 ;
      RECT 0.800 0.310 1.125 0.380 ;
      RECT 0.585 0.875 1.250 0.945 ;
      RECT 1.125 0.220 1.275 0.380 ;
      RECT 0.440 1.155 1.565 1.225 ;
      RECT 1.565 0.875 1.635 1.225 ;
      RECT 1.635 0.875 1.805 0.945 ;
      RECT 1.805 0.570 1.895 0.945 ;
  END
END INCLP3W111OF3X1

MACRO INCLP3W111OF3X2
  CLASS CORE ;
  FOREIGN INCLP3W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.675 0.590 0.810 0.805 ;
        RECT 0.810 0.735 1.910 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.870 1.370 0.945 ;
        RECT 1.370 0.870 1.600 1.180 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.585 1.530 0.670 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.700 0.870 1.975 1.155 ;
        RECT 1.975 0.150 2.045 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 0.995 0.340 1.485 ;
        RECT 0.340 1.315 1.655 1.485 ;
        RECT 1.655 1.220 1.885 1.485 ;
        RECT 1.885 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.335 0.250 ;
        RECT 0.335 -0.085 1.655 0.085 ;
        RECT 1.655 -0.085 1.885 0.385 ;
        RECT 1.885 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.135 1.235 ;
      RECT 0.135 0.655 0.340 0.930 ;
      RECT 0.200 0.315 0.405 0.590 ;
      RECT 0.405 0.315 0.475 1.080 ;
      RECT 0.540 0.450 0.610 0.895 ;
      RECT 0.400 0.175 1.105 0.250 ;
      RECT 0.445 1.145 1.105 1.225 ;
      RECT 0.475 0.315 1.170 0.385 ;
      RECT 0.475 1.010 1.170 1.080 ;
      RECT 1.170 0.225 1.305 0.385 ;
      RECT 1.170 1.010 1.305 1.250 ;
      RECT 0.610 0.450 1.655 0.520 ;
      RECT 1.655 0.450 1.910 0.670 ;
  END
END INCLP3W111OF3X2

MACRO INCLP3W111OF3X4
  CLASS CORE ;
  FOREIGN INCLP3W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.525 0.630 0.660 0.895 ;
        RECT 0.660 0.630 0.755 0.805 ;
        RECT 0.755 0.730 1.720 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.870 1.530 0.950 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046750 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.585 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105125 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.050 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.265 1.485 ;
        RECT 0.265 0.955 0.355 1.485 ;
        RECT 0.355 1.315 1.570 1.485 ;
        RECT 1.570 1.215 1.750 1.485 ;
        RECT 1.750 1.315 2.145 1.485 ;
        RECT 2.145 0.705 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.215 ;
        RECT 0.340 -0.085 1.565 0.085 ;
        RECT 1.565 -0.085 1.850 0.215 ;
        RECT 1.850 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.400 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.115 1.230 ;
      RECT 0.115 0.655 0.135 1.230 ;
      RECT 0.180 0.310 0.260 0.585 ;
      RECT 0.135 0.655 0.340 0.735 ;
      RECT 0.340 0.450 0.430 0.735 ;
      RECT 0.445 0.985 0.550 1.225 ;
      RECT 0.430 0.175 0.985 0.245 ;
      RECT 0.550 1.155 1.035 1.225 ;
      RECT 0.260 0.310 1.075 0.385 ;
      RECT 1.075 0.210 1.250 0.385 ;
      RECT 0.430 0.450 1.625 0.520 ;
      RECT 1.625 0.450 1.750 0.615 ;
      RECT 1.250 0.305 1.815 0.385 ;
      RECT 0.640 1.015 1.815 1.090 ;
      RECT 1.815 0.305 1.895 1.090 ;
  END
END INCLP3W111OF3X4

MACRO INCLP4W1111OF4X1
  CLASS CORE ;
  FOREIGN INCLP4W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.550 0.425 0.850 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.450 0.480 0.805 ;
        RECT 0.480 0.730 1.040 0.805 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.395 1.105 0.665 ;
        RECT 0.180 0.870 1.105 0.960 ;
        RECT 1.105 0.395 1.195 0.960 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.395 0.500 1.775 0.775 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.235 2.240 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.230 1.485 ;
        RECT 0.230 1.180 0.385 1.485 ;
        RECT 0.385 1.315 0.590 1.485 ;
        RECT 0.590 1.180 0.755 1.485 ;
        RECT 0.755 1.315 1.760 1.485 ;
        RECT 1.760 0.975 1.895 1.485 ;
        RECT 1.895 1.315 2.335 1.485 ;
        RECT 2.335 0.680 2.425 1.485 ;
        RECT 2.425 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.365 0.225 ;
        RECT 0.365 -0.085 0.590 0.085 ;
        RECT 0.590 -0.085 0.745 0.225 ;
        RECT 0.745 -0.085 1.795 0.085 ;
        RECT 1.795 -0.085 1.930 0.275 ;
        RECT 1.930 -0.085 2.335 0.085 ;
        RECT 2.335 -0.085 2.425 0.495 ;
        RECT 2.425 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.165 0.135 0.360 ;
      RECT 0.135 0.290 0.435 0.360 ;
      RECT 0.435 0.165 0.525 0.360 ;
      RECT 0.525 0.290 0.810 0.360 ;
      RECT 0.045 1.025 0.825 1.115 ;
      RECT 0.810 0.175 0.880 0.360 ;
      RECT 0.825 1.025 0.895 1.225 ;
      RECT 1.260 0.310 1.330 1.080 ;
      RECT 1.330 0.975 1.505 1.080 ;
      RECT 1.330 0.310 1.510 0.410 ;
      RECT 0.880 0.175 1.570 0.245 ;
      RECT 0.895 1.145 1.570 1.225 ;
      RECT 1.570 0.975 1.695 1.225 ;
      RECT 1.570 0.175 1.730 0.275 ;
      RECT 1.510 0.340 1.840 0.410 ;
      RECT 1.840 0.340 1.930 0.695 ;
      RECT 1.490 0.840 1.995 0.910 ;
      RECT 1.995 0.235 2.085 1.250 ;
  END
END INCLP4W1111OF4X1

MACRO INCLP4W1111OF4X2
  CLASS CORE ;
  FOREIGN INCLP4W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.350 0.595 0.650 0.810 ;
        RECT 0.650 0.595 0.835 0.685 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.325 0.435 0.900 0.525 ;
        RECT 0.900 0.435 1.025 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.260 0.965 ;
        RECT 0.260 0.875 1.090 0.965 ;
        RECT 1.090 0.535 1.180 0.965 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 1.380 0.535 1.465 0.875 ;
        RECT 1.465 0.805 1.580 0.875 ;
        RECT 1.580 0.805 1.715 1.015 ;
        RECT 1.715 0.805 1.815 0.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.805 2.335 1.105 ;
        RECT 2.335 0.195 2.425 1.105 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.225 0.355 1.485 ;
        RECT 0.355 1.315 0.580 1.485 ;
        RECT 0.580 1.225 0.780 1.485 ;
        RECT 0.780 1.315 1.780 1.485 ;
        RECT 1.780 0.940 1.915 1.485 ;
        RECT 1.915 1.315 2.150 1.485 ;
        RECT 2.150 1.170 2.265 1.485 ;
        RECT 2.265 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.170 ;
        RECT 0.355 -0.085 0.580 0.085 ;
        RECT 0.580 -0.085 0.780 0.170 ;
        RECT 0.780 -0.085 1.780 0.085 ;
        RECT 1.780 -0.085 1.915 0.335 ;
        RECT 1.915 -0.085 2.165 0.085 ;
        RECT 2.165 -0.085 2.265 0.400 ;
        RECT 2.265 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.140 0.305 ;
      RECT 0.045 1.080 0.140 1.250 ;
      RECT 0.140 0.235 0.425 0.305 ;
      RECT 0.425 0.150 0.515 0.305 ;
      RECT 1.245 0.370 1.315 1.015 ;
      RECT 1.315 0.370 1.515 0.470 ;
      RECT 1.315 0.940 1.515 1.015 ;
      RECT 0.515 0.235 1.575 0.305 ;
      RECT 1.530 0.535 1.670 0.740 ;
      RECT 1.575 0.235 1.715 0.335 ;
      RECT 0.140 1.080 1.715 1.160 ;
      RECT 1.515 0.400 1.810 0.470 ;
      RECT 1.810 0.400 1.915 0.595 ;
      RECT 1.670 0.660 1.995 0.740 ;
      RECT 1.995 0.300 2.085 1.180 ;
      RECT 2.085 0.300 2.100 0.730 ;
      RECT 2.100 0.465 2.265 0.730 ;
  END
END INCLP4W1111OF4X2

MACRO INCLP4W1111OF4X4
  CLASS CORE ;
  FOREIGN INCLP4W1111OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.430 0.770 0.635 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.360 0.725 0.895 0.805 ;
        RECT 0.895 0.455 1.005 0.805 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.135 0.730 0.270 0.950 ;
        RECT 0.270 0.870 1.095 0.950 ;
        RECT 1.095 0.645 1.185 0.950 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050750 ;
    PORT
      LAYER metal1 ;
        RECT 1.385 0.595 1.510 0.730 ;
        RECT 1.510 0.595 1.720 0.805 ;
        RECT 1.720 0.595 1.910 0.665 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105125 ;
    PORT
      LAYER metal1 ;
        RECT 2.340 0.230 2.430 1.080 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.240 0.375 1.485 ;
        RECT 0.375 1.315 0.585 1.485 ;
        RECT 0.585 1.240 0.805 1.485 ;
        RECT 0.805 1.315 1.810 1.485 ;
        RECT 1.810 1.035 1.905 1.485 ;
        RECT 1.905 1.315 2.160 1.485 ;
        RECT 2.160 0.725 2.250 1.485 ;
        RECT 2.250 1.315 2.525 1.485 ;
        RECT 2.525 0.725 2.615 1.485 ;
        RECT 2.615 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.170 ;
        RECT 0.340 -0.085 0.585 0.085 ;
        RECT 0.585 -0.085 0.805 0.170 ;
        RECT 0.805 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.905 0.365 ;
        RECT 1.905 -0.085 2.160 0.085 ;
        RECT 2.160 -0.085 2.250 0.410 ;
        RECT 2.250 -0.085 2.525 0.085 ;
        RECT 2.525 -0.085 2.615 0.440 ;
        RECT 2.615 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.340 ;
      RECT 0.125 0.260 0.430 0.340 ;
      RECT 0.430 0.175 0.510 0.340 ;
      RECT 0.510 0.260 0.895 0.340 ;
      RECT 0.895 0.175 0.975 0.340 ;
      RECT 1.250 0.310 1.320 0.950 ;
      RECT 1.320 0.310 1.515 0.390 ;
      RECT 0.975 0.175 1.605 0.245 ;
      RECT 1.605 0.175 1.695 0.365 ;
      RECT 0.045 1.040 1.720 1.175 ;
      RECT 1.320 0.870 1.810 0.950 ;
      RECT 1.810 0.730 1.910 0.950 ;
      RECT 1.510 0.455 1.995 0.530 ;
      RECT 1.995 0.310 2.000 0.530 ;
      RECT 2.000 0.310 2.075 1.175 ;
      RECT 2.075 0.500 2.250 0.635 ;
  END
END INCLP4W1111OF4X4

MACRO NCL1W1111OF4X1
  CLASS CORE ;
  FOREIGN NCL1W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.795 0.520 0.895 1.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.385 0.545 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.235 0.385 0.350 0.875 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.050 0.280 0.140 0.735 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 0.960 1.015 1.010 1.250 ;
        RECT 1.010 0.185 1.095 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.785 1.485 ;
        RECT 0.785 1.115 0.895 1.485 ;
        RECT 0.895 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.050 0.085 ;
        RECT 0.050 -0.085 0.170 0.215 ;
        RECT 0.170 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.545 0.185 ;
        RECT 0.545 -0.085 0.785 0.085 ;
        RECT 0.785 -0.085 0.895 0.255 ;
        RECT 0.895 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.050 0.940 0.200 1.215 ;
      RECT 0.235 0.160 0.325 0.320 ;
      RECT 0.325 0.250 0.615 0.320 ;
      RECT 0.615 0.160 0.635 0.320 ;
      RECT 0.200 0.940 0.635 1.010 ;
      RECT 0.635 0.160 0.705 1.010 ;
      RECT 0.705 0.320 0.935 0.455 ;
  END
END NCL1W1111OF4X1

MACRO NCL1W1111OF4X2
  CLASS CORE ;
  FOREIGN NCL1W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.385 0.785 0.595 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.660 0.760 1.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.230 0.385 0.510 1.015 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.050 0.280 0.140 0.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 1.005 0.170 1.095 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.770 1.485 ;
        RECT 0.770 1.215 0.940 1.485 ;
        RECT 0.940 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.055 0.085 ;
        RECT 0.055 -0.085 0.185 0.215 ;
        RECT 0.185 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.545 0.180 ;
        RECT 0.545 -0.085 0.770 0.085 ;
        RECT 0.770 -0.085 0.940 0.185 ;
        RECT 0.940 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.940 0.135 1.250 ;
      RECT 0.135 1.080 0.185 1.250 ;
      RECT 0.250 0.165 0.335 0.320 ;
      RECT 0.335 0.250 0.615 0.320 ;
      RECT 0.615 0.165 0.705 0.320 ;
      RECT 0.705 0.250 0.850 0.320 ;
      RECT 0.185 1.080 0.850 1.150 ;
      RECT 0.850 0.250 0.940 1.150 ;
  END
END NCL1W1111OF4X2

MACRO NCL1W111OF3X1
  CLASS CORE ;
  FOREIGN NCL1W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.385 0.785 0.920 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.350 0.385 0.510 0.920 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021000 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.385 0.260 0.875 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.042350 ;
    PORT
      LAYER metal1 ;
        RECT 1.010 0.150 1.095 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.660 1.485 ;
        RECT 0.660 1.120 0.750 1.485 ;
        RECT 0.750 1.120 0.945 1.225 ;
        RECT 0.750 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.260 0.085 ;
        RECT 0.260 -0.085 0.395 0.185 ;
        RECT 0.395 -0.085 0.800 0.085 ;
        RECT 0.800 -0.085 0.945 0.185 ;
        RECT 0.945 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.055 0.150 0.195 0.320 ;
      RECT 0.055 0.985 0.350 1.250 ;
      RECT 0.195 0.250 0.460 0.320 ;
      RECT 0.460 0.150 0.735 0.320 ;
      RECT 0.735 0.250 0.875 0.320 ;
      RECT 0.350 0.985 0.875 1.055 ;
      RECT 0.875 0.250 0.945 1.055 ;
  END
END NCL1W111OF3X1

MACRO NCL1W111OF3X2
  CLASS CORE ;
  FOREIGN NCL1W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021750 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.385 0.780 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021750 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.385 0.540 0.875 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021750 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.350 0.875 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.005 0.155 1.095 1.240 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.750 1.485 ;
        RECT 0.750 1.110 0.940 1.485 ;
        RECT 0.940 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.385 0.085 ;
        RECT 0.385 -0.085 0.520 0.185 ;
        RECT 0.520 -0.085 0.795 0.085 ;
        RECT 0.795 -0.085 0.940 0.185 ;
        RECT 0.940 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.155 0.320 0.320 ;
      RECT 0.045 0.940 0.370 1.150 ;
      RECT 0.320 0.250 0.590 0.320 ;
      RECT 0.590 0.155 0.725 0.320 ;
      RECT 0.725 0.250 0.870 0.320 ;
      RECT 0.370 0.940 0.870 1.040 ;
      RECT 0.870 0.250 0.940 1.040 ;
  END
END NCL1W111OF3X2

MACRO NCL1W111OF3X4
  CLASS CORE ;
  FOREIGN NCL1W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.455 0.595 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.735 0.440 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.095 0.455 0.270 0.660 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105850 ;
    PORT
      LAYER metal1 ;
        RECT 0.820 0.215 0.910 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.550 1.485 ;
        RECT 0.550 1.195 0.720 1.485 ;
        RECT 0.720 1.315 1.005 1.485 ;
        RECT 1.005 0.815 1.095 1.485 ;
        RECT 1.095 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.210 0.085 ;
        RECT 0.210 -0.085 0.345 0.225 ;
        RECT 0.345 -0.085 0.605 0.085 ;
        RECT 0.605 -0.085 0.740 0.225 ;
        RECT 0.740 -0.085 1.005 0.085 ;
        RECT 1.005 -0.085 1.095 0.445 ;
        RECT 1.095 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.935 0.115 1.225 ;
      RECT 0.045 0.175 0.125 0.390 ;
      RECT 0.115 1.025 0.145 1.225 ;
      RECT 0.125 0.310 0.435 0.390 ;
      RECT 0.435 0.175 0.515 0.390 ;
      RECT 0.515 0.310 0.665 0.390 ;
      RECT 0.145 1.025 0.665 1.105 ;
      RECT 0.665 0.310 0.745 1.105 ;
  END
END NCL1W111OF3X4

MACRO NCL1W11OF2X1
  CLASS CORE ;
  FOREIGN NCL1W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019250 ;
    PORT
      LAYER metal1 ;
        RECT 0.050 0.375 0.140 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019250 ;
    PORT
      LAYER metal1 ;
        RECT 0.240 0.385 0.405 0.875 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.150 0.715 1.240 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.355 1.485 ;
        RECT 0.355 1.115 0.565 1.485 ;
        RECT 0.565 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.140 0.310 ;
        RECT 0.140 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.565 0.185 ;
        RECT 0.565 -0.085 0.760 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.940 0.140 1.240 ;
      RECT 0.240 0.150 0.330 0.320 ;
      RECT 0.330 0.250 0.495 0.320 ;
      RECT 0.140 0.940 0.495 1.035 ;
      RECT 0.495 0.250 0.565 1.035 ;
  END
END NCL1W11OF2X1

MACRO NCL1W11OF2X2
  CLASS CORE ;
  FOREIGN NCL1W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.320 0.135 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019250 ;
    PORT
      LAYER metal1 ;
        RECT 0.240 0.385 0.405 0.735 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.081400 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.155 0.715 1.240 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.405 1.485 ;
        RECT 0.405 0.940 0.565 1.485 ;
        RECT 0.565 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.255 ;
        RECT 0.135 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.565 0.185 ;
        RECT 0.565 -0.085 0.760 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.800 0.135 1.100 ;
      RECT 0.225 0.155 0.315 0.320 ;
      RECT 0.315 0.250 0.495 0.320 ;
      RECT 0.135 0.800 0.495 0.870 ;
      RECT 0.495 0.250 0.565 0.870 ;
  END
END NCL1W11OF2X2

MACRO NCL1W11OF2X4
  CLASS CORE ;
  FOREIGN NCL1W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.370 0.135 0.645 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020250 ;
    PORT
      LAYER metal1 ;
        RECT 0.240 0.385 0.405 0.875 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.106575 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.175 0.720 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.410 1.485 ;
        RECT 0.410 1.080 0.545 1.485 ;
        RECT 0.545 1.315 0.810 1.485 ;
        RECT 0.810 0.845 0.900 1.485 ;
        RECT 0.900 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.280 ;
        RECT 0.135 -0.085 0.410 0.085 ;
        RECT 0.410 -0.085 0.545 0.180 ;
        RECT 0.545 -0.085 0.810 0.085 ;
        RECT 0.810 -0.085 0.900 0.445 ;
        RECT 0.900 -0.085 0.950 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.820 0.150 1.110 ;
      RECT 0.150 0.940 0.155 1.110 ;
      RECT 0.235 0.170 0.320 0.320 ;
      RECT 0.320 0.245 0.495 0.320 ;
      RECT 0.155 0.940 0.495 1.015 ;
      RECT 0.495 0.245 0.565 1.015 ;
  END
END NCL1W11OF2X4

MACRO NCL1W1OF1X1
  CLASS CORE ;
  FOREIGN NCL1W1OF1X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.018000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.385 0.195 0.875 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.160 0.510 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.075 0.355 1.485 ;
        RECT 0.355 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.185 ;
        RECT 0.355 -0.085 0.570 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.160 0.135 0.320 ;
      RECT 0.045 0.940 0.135 1.100 ;
      RECT 0.135 0.250 0.285 0.320 ;
      RECT 0.135 0.940 0.285 1.010 ;
      RECT 0.285 0.250 0.355 1.010 ;
  END
END NCL1W1OF1X1

MACRO NCL1W1OF1X2
  CLASS CORE ;
  FOREIGN NCL1W1OF1X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.570 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019000 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.380 0.190 0.735 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080850 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.155 0.510 1.175 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 0.945 0.355 1.485 ;
        RECT 0.355 1.315 0.570 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.175 ;
        RECT 0.355 -0.085 0.570 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.155 0.135 0.315 ;
      RECT 0.045 0.805 0.135 1.175 ;
      RECT 0.135 0.245 0.285 0.315 ;
      RECT 0.135 0.805 0.285 0.875 ;
      RECT 0.285 0.245 0.355 0.875 ;
  END
END NCL1W1OF1X2

MACRO NCL1W1OF1X4
  CLASS CORE ;
  FOREIGN NCL1W1OF1X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.018000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.195 1.015 ;
    END
  END A
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105125 ;
    PORT
      LAYER metal1 ;
        RECT 0.420 0.165 0.510 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 1.215 0.355 1.485 ;
        RECT 0.355 1.315 0.600 1.485 ;
        RECT 0.600 0.870 0.695 1.485 ;
        RECT 0.695 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.290 ;
        RECT 0.355 -0.085 0.600 0.085 ;
        RECT 0.600 -0.085 0.695 0.455 ;
        RECT 0.695 -0.085 0.760 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.165 0.135 0.460 ;
      RECT 0.045 1.080 0.135 1.250 ;
      RECT 0.135 0.390 0.285 0.460 ;
      RECT 0.135 1.080 0.285 1.150 ;
      RECT 0.285 0.390 0.355 1.150 ;
  END
END NCL1W1OF1X4

MACRO NCL2W11OF2X1
  CLASS CORE ;
  FOREIGN NCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.041750 ;
    PORT
      LAYER metal1 ;
        RECT 0.170 0.805 0.710 1.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.041750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.510 0.960 0.715 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 1.360 0.385 1.575 0.685 ;
        RECT 1.575 0.155 1.665 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.065 0.125 1.485 ;
        RECT 0.125 1.315 0.395 1.485 ;
        RECT 0.395 1.240 0.540 1.485 ;
        RECT 0.540 1.315 1.380 1.485 ;
        RECT 1.380 0.820 1.470 1.485 ;
        RECT 1.470 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.050 0.085 ;
        RECT 0.050 -0.085 0.140 0.400 ;
        RECT 0.140 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.540 0.280 ;
        RECT 0.540 -0.085 1.360 0.085 ;
        RECT 1.360 -0.085 1.470 0.310 ;
        RECT 1.470 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.255 0.310 0.415 ;
      RECT 0.205 1.105 0.605 1.175 ;
      RECT 0.310 0.345 0.640 0.415 ;
      RECT 0.605 1.105 0.675 1.225 ;
      RECT 0.640 0.175 0.710 0.415 ;
      RECT 0.780 0.310 0.940 0.445 ;
      RECT 0.780 0.780 0.940 1.070 ;
      RECT 0.710 0.175 1.005 0.245 ;
      RECT 0.675 1.155 1.005 1.225 ;
      RECT 0.940 0.375 1.050 0.445 ;
      RECT 0.940 0.780 1.050 0.955 ;
      RECT 1.005 0.175 1.140 0.310 ;
      RECT 1.050 0.375 1.140 0.955 ;
      RECT 1.005 1.020 1.140 1.225 ;
      RECT 1.205 0.155 1.295 1.225 ;
  END
END NCL2W11OF2X1

MACRO NCL2W11OF2X2
  CLASS CORE ;
  FOREIGN NCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.730 0.820 0.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.575 0.995 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.520 0.440 1.765 0.740 ;
        RECT 1.765 0.245 1.855 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.055 1.485 ;
        RECT 0.055 0.885 0.150 1.485 ;
        RECT 0.150 1.315 0.400 1.485 ;
        RECT 0.400 1.040 0.685 1.485 ;
        RECT 0.685 1.315 1.520 1.485 ;
        RECT 1.520 0.885 1.660 1.485 ;
        RECT 1.660 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.070 0.085 ;
        RECT 0.070 -0.085 0.180 0.430 ;
        RECT 0.180 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.595 0.370 ;
        RECT 0.595 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.660 0.365 ;
        RECT 1.660 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.245 0.300 0.360 0.510 ;
      RECT 0.360 0.440 0.660 0.510 ;
      RECT 0.660 0.175 0.735 0.510 ;
      RECT 0.215 0.885 0.750 0.975 ;
      RECT 0.750 0.885 0.820 1.225 ;
      RECT 0.805 0.335 1.060 0.510 ;
      RECT 0.885 0.730 1.060 1.090 ;
      RECT 1.060 0.335 1.100 1.090 ;
      RECT 1.100 0.335 1.130 0.855 ;
      RECT 0.820 1.155 1.165 1.225 ;
      RECT 0.735 0.175 1.195 0.245 ;
      RECT 1.195 0.175 1.300 0.430 ;
      RECT 1.130 0.555 1.300 0.855 ;
      RECT 1.165 0.920 1.300 1.225 ;
      RECT 1.365 0.245 1.455 1.155 ;
  END
END NCL2W11OF2X2

MACRO NCL2W11OF2X4
  CLASS CORE ;
  FOREIGN NCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.735 0.370 0.825 ;
        RECT 0.370 0.735 0.590 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.330 0.455 0.805 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.565 0.175 1.660 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.970 0.125 1.485 ;
        RECT 0.125 1.315 0.395 1.485 ;
        RECT 0.395 1.160 0.535 1.485 ;
        RECT 0.535 1.315 1.385 1.485 ;
        RECT 1.385 0.745 1.475 1.485 ;
        RECT 1.475 1.315 1.765 1.485 ;
        RECT 1.765 0.675 1.855 1.485 ;
        RECT 1.855 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.305 ;
        RECT 0.135 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.530 0.195 ;
        RECT 0.530 -0.085 1.385 0.085 ;
        RECT 1.385 -0.085 1.475 0.455 ;
        RECT 1.475 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.855 0.445 ;
        RECT 1.855 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.195 0.305 0.365 ;
      RECT 0.205 1.010 0.305 1.250 ;
      RECT 0.305 0.285 0.620 0.365 ;
      RECT 0.305 1.010 0.625 1.090 ;
      RECT 0.620 0.175 0.700 0.365 ;
      RECT 0.625 1.010 0.705 1.225 ;
      RECT 0.790 0.310 0.870 0.390 ;
      RECT 0.795 0.755 0.870 1.055 ;
      RECT 0.870 0.310 0.950 1.055 ;
      RECT 0.700 0.175 1.035 0.245 ;
      RECT 0.705 1.145 1.040 1.225 ;
      RECT 1.035 0.175 1.115 0.335 ;
      RECT 0.950 0.440 1.125 0.575 ;
      RECT 1.030 0.665 1.205 0.870 ;
      RECT 1.040 0.950 1.245 1.225 ;
      RECT 1.205 0.315 1.295 0.870 ;
  END
END NCL2W11OF2X4

MACRO NCL2W211OF3X1
  CLASS CORE ;
  FOREIGN NCL2W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024250 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.595 1.595 0.675 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.510 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.110 0.825 0.600 0.915 ;
        RECT 0.600 0.525 0.890 0.915 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.385 1.955 0.595 ;
        RECT 1.955 0.175 2.045 0.960 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.005 0.125 1.485 ;
        RECT 0.125 1.315 0.405 1.485 ;
        RECT 0.405 1.180 0.540 1.485 ;
        RECT 0.540 1.315 1.770 1.485 ;
        RECT 1.770 0.685 1.860 1.485 ;
        RECT 1.860 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.300 ;
        RECT 0.135 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.540 0.265 ;
        RECT 0.540 -0.085 1.365 0.085 ;
        RECT 1.365 -0.085 1.455 0.215 ;
        RECT 1.455 -0.085 1.770 0.085 ;
        RECT 1.770 -0.085 1.860 0.295 ;
        RECT 1.860 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.225 0.315 0.435 ;
      RECT 0.315 0.355 0.630 0.435 ;
      RECT 0.630 0.175 0.710 0.435 ;
      RECT 0.800 0.315 0.980 0.435 ;
      RECT 0.980 0.315 1.060 0.955 ;
      RECT 0.215 1.020 1.080 1.090 ;
      RECT 0.710 0.175 1.095 0.250 ;
      RECT 1.060 0.875 1.170 0.955 ;
      RECT 1.060 0.315 1.185 0.395 ;
      RECT 1.150 0.460 1.230 0.810 ;
      RECT 1.170 0.875 1.230 1.065 ;
      RECT 1.185 0.175 1.275 0.395 ;
      RECT 0.725 1.155 1.290 1.225 ;
      RECT 1.230 0.900 1.485 1.065 ;
      RECT 1.275 0.305 1.525 0.395 ;
      RECT 1.230 0.460 1.590 0.530 ;
      RECT 1.230 0.740 1.665 0.810 ;
      RECT 1.590 0.175 1.680 0.530 ;
  END
END NCL2W211OF3X1

MACRO NCL2W211OF3X2
  CLASS CORE ;
  FOREIGN NCL2W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.455 1.355 0.590 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.510 0.760 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.855 0.600 0.945 ;
        RECT 0.600 0.525 0.815 0.945 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078100 ;
    PORT
      LAYER metal1 ;
        RECT 1.775 0.435 1.955 0.525 ;
        RECT 1.955 0.215 2.045 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.130 1.485 ;
        RECT 0.130 1.315 0.450 1.485 ;
        RECT 0.450 1.180 0.550 1.485 ;
        RECT 0.550 1.315 1.775 1.485 ;
        RECT 1.775 0.615 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.300 ;
        RECT 0.135 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.265 ;
        RECT 0.550 -0.085 1.360 0.085 ;
        RECT 1.360 -0.085 1.495 0.220 ;
        RECT 1.495 -0.085 1.775 0.085 ;
        RECT 1.775 -0.085 1.865 0.300 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.215 0.325 0.435 ;
      RECT 0.220 1.020 0.360 1.225 ;
      RECT 0.325 0.355 0.630 0.435 ;
      RECT 0.630 0.175 0.710 0.435 ;
      RECT 0.800 0.315 0.905 0.405 ;
      RECT 0.905 0.315 0.985 0.930 ;
      RECT 0.710 0.175 1.090 0.250 ;
      RECT 0.360 1.020 1.090 1.090 ;
      RECT 0.985 0.315 1.180 0.390 ;
      RECT 1.180 0.215 1.270 0.390 ;
      RECT 0.745 1.155 1.285 1.225 ;
      RECT 1.270 0.310 1.445 0.390 ;
      RECT 0.985 0.850 1.480 0.930 ;
      RECT 1.445 0.310 1.525 0.490 ;
      RECT 1.075 0.680 1.590 0.760 ;
      RECT 1.590 0.215 1.685 0.760 ;
      RECT 1.480 0.850 1.685 1.210 ;
  END
END NCL2W211OF3X2

MACRO NCL2W211OF3X4
  CLASS CORE ;
  FOREIGN NCL2W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.315 1.530 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.510 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.855 0.600 0.945 ;
        RECT 0.600 0.635 0.850 0.945 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.955 0.245 2.045 1.090 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.130 1.485 ;
        RECT 0.130 1.315 0.450 1.485 ;
        RECT 0.450 1.180 0.625 1.485 ;
        RECT 0.625 1.315 1.775 1.485 ;
        RECT 1.775 0.675 1.865 1.485 ;
        RECT 1.865 1.315 2.145 1.485 ;
        RECT 2.145 0.705 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.305 ;
        RECT 0.130 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.560 0.265 ;
        RECT 0.560 -0.085 1.345 0.085 ;
        RECT 1.345 -0.085 1.620 0.225 ;
        RECT 1.620 -0.085 1.775 0.085 ;
        RECT 1.775 -0.085 1.865 0.485 ;
        RECT 1.865 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.465 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.265 0.310 0.435 ;
      RECT 0.220 1.020 0.360 1.225 ;
      RECT 0.310 0.355 0.650 0.435 ;
      RECT 0.650 0.175 0.730 0.435 ;
      RECT 0.825 0.345 0.915 0.545 ;
      RECT 0.915 0.465 0.940 0.545 ;
      RECT 0.730 0.175 1.005 0.255 ;
      RECT 0.940 0.465 1.020 0.955 ;
      RECT 1.005 0.175 1.095 0.375 ;
      RECT 0.360 1.020 1.135 1.090 ;
      RECT 1.020 0.465 1.175 0.545 ;
      RECT 1.175 0.195 1.255 0.545 ;
      RECT 0.800 1.155 1.285 1.225 ;
      RECT 1.020 0.875 1.375 0.955 ;
      RECT 1.110 0.730 1.595 0.810 ;
      RECT 1.375 0.875 1.650 1.225 ;
      RECT 1.595 0.400 1.685 0.810 ;
  END
END NCL2W211OF3X4

MACRO NCL3W111OF3X1
  CLASS CORE ;
  FOREIGN NCL3W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.590 0.595 0.700 0.875 ;
        RECT 0.700 0.595 1.320 0.665 ;
        RECT 1.320 0.445 1.570 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048000 ;
    PORT
      LAYER metal1 ;
        RECT 0.935 0.730 1.150 0.945 ;
        RECT 1.150 0.855 1.265 0.945 ;
        RECT 1.265 0.730 1.530 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.445 1.255 0.530 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.042350 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.150 1.855 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.200 1.485 ;
        RECT 0.200 0.970 0.325 1.485 ;
        RECT 0.325 1.315 1.520 1.485 ;
        RECT 1.520 1.145 1.705 1.485 ;
        RECT 1.705 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.235 0.085 ;
        RECT 0.235 -0.085 0.345 0.330 ;
        RECT 0.345 -0.085 1.560 0.085 ;
        RECT 1.560 -0.085 1.705 0.245 ;
        RECT 1.705 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.275 0.135 0.465 ;
      RECT 0.045 0.835 0.135 1.250 ;
      RECT 0.115 0.530 0.215 0.770 ;
      RECT 0.135 0.395 0.280 0.465 ;
      RECT 0.135 0.835 0.390 0.905 ;
      RECT 0.280 0.395 0.440 0.635 ;
      RECT 0.215 0.700 0.455 0.770 ;
      RECT 0.425 0.175 0.515 0.330 ;
      RECT 0.455 0.700 0.525 1.080 ;
      RECT 0.525 1.010 0.750 1.080 ;
      RECT 0.750 0.920 0.840 1.080 ;
      RECT 0.515 0.175 0.920 0.245 ;
      RECT 0.390 1.145 0.945 1.225 ;
      RECT 0.580 0.310 0.985 0.380 ;
      RECT 0.840 1.010 1.010 1.080 ;
      RECT 1.010 1.010 1.125 1.250 ;
      RECT 0.985 0.220 1.495 0.380 ;
      RECT 1.495 0.310 1.635 0.380 ;
      RECT 1.125 1.010 1.635 1.080 ;
      RECT 1.635 0.310 1.705 1.080 ;
  END
END NCL3W111OF3X1

MACRO NCL3W111OF3X2
  CLASS CORE ;
  FOREIGN NCL3W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.730 1.405 0.805 ;
        RECT 1.405 0.505 1.570 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.870 1.540 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.575 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.150 1.855 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.190 1.485 ;
        RECT 0.190 1.145 0.335 1.485 ;
        RECT 0.335 1.315 1.520 1.485 ;
        RECT 1.520 1.165 1.705 1.485 ;
        RECT 1.705 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.360 0.340 ;
        RECT 0.360 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.705 0.260 ;
        RECT 1.705 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.290 0.125 1.145 ;
      RECT 0.125 0.290 0.135 0.650 ;
      RECT 0.190 0.715 0.280 1.080 ;
      RECT 0.135 0.445 0.475 0.650 ;
      RECT 0.425 0.185 0.525 0.340 ;
      RECT 0.590 0.325 0.765 0.485 ;
      RECT 0.525 0.185 0.830 0.255 ;
      RECT 0.830 0.185 0.925 0.340 ;
      RECT 0.400 1.145 0.945 1.225 ;
      RECT 0.765 0.415 0.990 0.485 ;
      RECT 0.280 1.010 1.010 1.080 ;
      RECT 1.010 1.010 1.130 1.250 ;
      RECT 0.990 0.325 1.150 0.485 ;
      RECT 1.150 0.325 1.635 0.395 ;
      RECT 1.130 1.010 1.635 1.100 ;
      RECT 1.635 0.325 1.705 1.100 ;
  END
END NCL3W111OF3X2

MACRO NCL3W111OF3X4
  CLASS CORE ;
  FOREIGN NCL3W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.540 0.730 1.465 0.805 ;
        RECT 1.465 0.465 1.555 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.870 0.870 1.465 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.745 0.585 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.107300 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.170 1.860 1.235 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.220 1.485 ;
        RECT 0.220 0.960 0.300 1.485 ;
        RECT 0.300 1.315 1.520 1.485 ;
        RECT 1.520 1.205 1.680 1.485 ;
        RECT 1.680 1.315 1.955 1.485 ;
        RECT 1.955 0.890 2.045 1.485 ;
        RECT 2.045 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.220 0.085 ;
        RECT 0.220 -0.085 0.310 0.355 ;
        RECT 0.310 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.660 0.205 ;
        RECT 1.660 -0.085 1.955 0.085 ;
        RECT 1.955 -0.085 2.045 0.355 ;
        RECT 2.045 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.295 0.130 0.530 ;
      RECT 0.045 0.740 0.130 1.235 ;
      RECT 0.130 0.740 0.335 0.875 ;
      RECT 0.135 0.595 0.400 0.675 ;
      RECT 0.130 0.445 0.435 0.530 ;
      RECT 0.400 0.595 0.475 1.080 ;
      RECT 0.400 0.175 0.490 0.355 ;
      RECT 0.580 0.345 0.725 0.500 ;
      RECT 0.490 0.175 0.815 0.255 ;
      RECT 0.390 1.145 0.905 1.225 ;
      RECT 0.815 0.175 0.920 0.330 ;
      RECT 0.475 1.010 0.995 1.080 ;
      RECT 0.725 0.420 1.010 0.500 ;
      RECT 0.995 1.010 1.125 1.250 ;
      RECT 1.010 0.295 1.155 0.500 ;
      RECT 1.155 0.295 1.620 0.375 ;
      RECT 1.125 1.035 1.620 1.115 ;
      RECT 1.620 0.295 1.700 1.115 ;
  END
END NCL3W111OF3X4

MACRO NCL3W211OF3X1
  CLASS CORE ;
  FOREIGN NCL3W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.455 0.580 0.710 ;
        RECT 0.580 0.640 1.135 0.710 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.505 0.775 1.130 0.845 ;
        RECT 1.130 0.775 1.200 0.945 ;
        RECT 1.200 0.665 1.340 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 0.090 0.805 0.390 0.980 ;
        RECT 0.390 0.910 0.825 0.980 ;
        RECT 0.825 0.910 0.895 1.225 ;
        RECT 0.895 1.155 1.590 1.225 ;
        RECT 1.590 0.880 1.690 1.225 ;
        RECT 1.690 0.880 1.870 0.970 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.235 2.235 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.270 1.485 ;
        RECT 0.270 1.205 0.390 1.485 ;
        RECT 0.390 1.315 1.780 1.485 ;
        RECT 1.780 1.060 1.870 1.485 ;
        RECT 1.870 1.315 1.965 1.485 ;
        RECT 1.965 0.640 2.055 1.485 ;
        RECT 2.055 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.080 0.085 ;
        RECT 0.080 -0.085 0.180 0.205 ;
        RECT 0.180 -0.085 0.455 0.085 ;
        RECT 0.455 -0.085 0.545 0.205 ;
        RECT 0.545 -0.085 1.365 0.085 ;
        RECT 1.365 -0.085 1.505 0.170 ;
        RECT 1.505 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.055 0.480 ;
        RECT 2.055 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 1.045 0.180 1.250 ;
      RECT 0.270 0.175 0.365 0.365 ;
      RECT 0.180 1.045 0.620 1.115 ;
      RECT 0.365 0.295 0.635 0.365 ;
      RECT 0.635 0.175 0.725 0.365 ;
      RECT 0.620 1.045 0.760 1.250 ;
      RECT 0.790 0.175 0.860 0.575 ;
      RECT 0.860 0.175 1.095 0.280 ;
      RECT 1.185 0.170 1.275 0.305 ;
      RECT 0.860 0.505 1.430 0.575 ;
      RECT 0.980 1.010 1.430 1.080 ;
      RECT 1.430 0.505 1.500 1.080 ;
      RECT 1.275 0.235 1.595 0.305 ;
      RECT 1.500 0.505 1.700 0.775 ;
      RECT 0.945 0.370 1.765 0.440 ;
      RECT 1.595 0.175 1.870 0.305 ;
      RECT 1.765 0.370 1.870 0.790 ;
  END
END NCL3W211OF3X1

MACRO NCL3W211OF3X2
  CLASS CORE ;
  FOREIGN NCL3W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.400 0.580 0.640 ;
        RECT 0.580 0.400 0.710 0.750 ;
        RECT 0.710 0.660 1.130 0.750 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.580 0.815 1.200 0.905 ;
        RECT 1.200 0.630 1.345 0.905 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.230 0.705 0.510 1.040 ;
        RECT 0.510 0.970 0.815 1.040 ;
        RECT 0.815 0.970 0.885 1.225 ;
        RECT 0.885 1.155 1.545 1.225 ;
        RECT 1.545 0.715 1.615 1.225 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.077000 ;
    PORT
      LAYER metal1 ;
        RECT 1.925 0.360 2.145 0.630 ;
        RECT 2.145 0.225 2.235 1.170 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.230 1.485 ;
        RECT 0.230 1.240 0.375 1.485 ;
        RECT 0.375 1.315 1.680 1.485 ;
        RECT 1.680 0.990 1.885 1.485 ;
        RECT 1.885 1.315 1.975 1.485 ;
        RECT 1.975 0.700 2.065 1.485 ;
        RECT 2.065 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.075 0.085 ;
        RECT 0.075 -0.085 0.165 0.215 ;
        RECT 0.165 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.560 0.175 ;
        RECT 0.560 -0.085 1.330 0.085 ;
        RECT 1.330 -0.085 1.485 0.160 ;
        RECT 1.485 -0.085 1.925 0.085 ;
        RECT 1.925 -0.085 2.065 0.295 ;
        RECT 2.065 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.230 0.150 0.335 0.310 ;
      RECT 0.335 0.240 0.625 0.310 ;
      RECT 0.625 0.150 0.715 0.310 ;
      RECT 0.045 1.105 0.750 1.175 ;
      RECT 0.780 0.150 0.850 0.565 ;
      RECT 0.850 0.150 1.060 0.295 ;
      RECT 1.160 0.150 1.260 0.295 ;
      RECT 0.850 0.495 1.410 0.565 ;
      RECT 0.950 1.000 1.410 1.090 ;
      RECT 1.410 0.495 1.480 1.090 ;
      RECT 1.260 0.225 1.550 0.295 ;
      RECT 1.550 0.150 1.680 0.295 ;
      RECT 1.480 0.495 1.700 0.645 ;
      RECT 0.915 0.360 1.765 0.430 ;
      RECT 1.765 0.225 1.855 0.920 ;
  END
END NCL3W211OF3X2

MACRO NCL3W211OF3X4
  CLASS CORE ;
  FOREIGN NCL3W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.160 0.430 0.575 0.635 ;
        RECT 0.575 0.430 0.750 0.775 ;
        RECT 0.750 0.695 1.145 0.775 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.545 0.865 1.235 0.945 ;
        RECT 1.235 0.670 1.390 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.250 0.725 0.455 1.085 ;
        RECT 0.455 1.010 0.840 1.085 ;
        RECT 0.840 1.010 0.920 1.225 ;
        RECT 0.920 1.155 1.615 1.225 ;
        RECT 1.615 0.780 1.695 1.225 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.245 2.235 1.085 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.235 1.485 ;
        RECT 0.235 1.290 0.400 1.485 ;
        RECT 0.400 1.315 1.785 1.485 ;
        RECT 1.785 1.035 1.875 1.485 ;
        RECT 1.875 1.315 1.965 1.485 ;
        RECT 1.965 0.670 2.055 1.485 ;
        RECT 2.055 1.315 2.335 1.485 ;
        RECT 2.335 0.725 2.425 1.485 ;
        RECT 2.425 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.160 0.215 ;
        RECT 0.160 -0.085 0.440 0.085 ;
        RECT 0.440 -0.085 0.575 0.170 ;
        RECT 0.575 -0.085 1.380 0.085 ;
        RECT 1.380 -0.085 1.525 0.160 ;
        RECT 1.525 -0.085 1.965 0.085 ;
        RECT 1.965 -0.085 2.055 0.470 ;
        RECT 2.055 -0.085 2.335 0.085 ;
        RECT 2.335 -0.085 2.425 0.470 ;
        RECT 2.425 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.950 0.160 1.225 ;
      RECT 0.260 0.175 0.350 0.340 ;
      RECT 0.350 0.260 0.665 0.340 ;
      RECT 0.665 0.175 0.750 0.340 ;
      RECT 0.160 1.150 0.770 1.225 ;
      RECT 0.840 0.175 0.930 0.605 ;
      RECT 0.995 0.305 1.085 0.470 ;
      RECT 1.195 0.175 1.290 0.330 ;
      RECT 0.930 0.535 1.455 0.605 ;
      RECT 0.995 1.010 1.455 1.090 ;
      RECT 1.455 0.535 1.535 1.090 ;
      RECT 1.290 0.250 1.615 0.330 ;
      RECT 1.535 0.535 1.720 0.680 ;
      RECT 1.085 0.395 1.785 0.470 ;
      RECT 1.615 0.175 1.825 0.330 ;
      RECT 1.785 0.395 1.875 0.945 ;
  END
END NCL3W211OF3X4

MACRO NCL3W3111OF4X1
  CLASS CORE ;
  FOREIGN NCL3W3111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.650 0.135 0.945 ;
        RECT 0.135 0.875 0.370 0.945 ;
        RECT 0.370 0.875 0.770 1.225 ;
        RECT 0.770 0.875 1.510 0.945 ;
        RECT 1.510 0.730 1.720 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 0.295 0.595 1.340 0.665 ;
        RECT 1.340 0.460 1.570 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 0.470 0.730 1.340 0.810 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.455 0.825 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.044975 ;
    PORT
      LAYER metal1 ;
        RECT 2.305 0.500 2.525 0.590 ;
        RECT 2.525 0.245 2.615 1.015 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.010 0.135 1.485 ;
        RECT 0.135 1.315 1.920 1.485 ;
        RECT 1.920 1.010 2.055 1.485 ;
        RECT 2.055 1.315 2.305 1.485 ;
        RECT 2.305 0.655 2.420 1.485 ;
        RECT 2.420 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.355 0.255 ;
        RECT 0.355 -0.085 1.925 0.085 ;
        RECT 1.925 -0.085 2.055 0.335 ;
        RECT 2.055 -0.085 2.305 0.085 ;
        RECT 2.305 -0.085 2.420 0.435 ;
        RECT 2.420 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.230 0.135 0.390 ;
      RECT 0.135 0.320 0.685 0.390 ;
      RECT 0.685 0.215 0.795 0.390 ;
      RECT 0.795 0.305 0.855 0.390 ;
      RECT 0.855 0.305 0.885 0.395 ;
      RECT 0.935 0.175 1.070 0.260 ;
      RECT 0.885 0.325 1.115 0.395 ;
      RECT 1.115 0.310 1.635 0.395 ;
      RECT 1.115 1.145 1.655 1.225 ;
      RECT 1.635 0.310 1.705 0.625 ;
      RECT 1.070 0.175 1.770 0.245 ;
      RECT 1.705 0.490 1.785 0.625 ;
      RECT 0.895 1.010 1.785 1.080 ;
      RECT 1.785 0.490 1.855 1.080 ;
      RECT 1.770 0.175 1.860 0.335 ;
      RECT 1.855 0.490 2.095 0.625 ;
      RECT 1.920 0.690 2.160 0.945 ;
      RECT 2.160 0.320 2.240 0.945 ;
  END
END NCL3W3111OF4X1

MACRO NCL3W3111OF4X2
  CLASS CORE ;
  FOREIGN NCL3W3111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.660 0.225 0.945 ;
        RECT 0.225 0.875 0.440 0.945 ;
        RECT 0.440 0.875 0.740 1.165 ;
        RECT 0.740 0.875 1.580 0.945 ;
        RECT 1.580 0.665 1.720 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051250 ;
    PORT
      LAYER metal1 ;
        RECT 0.290 0.595 1.320 0.665 ;
        RECT 1.320 0.455 1.515 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051250 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.730 1.390 0.810 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051250 ;
    PORT
      LAYER metal1 ;
        RECT 0.550 0.445 0.960 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079750 ;
    PORT
      LAYER metal1 ;
        RECT 2.525 0.245 2.615 1.165 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.010 0.135 1.485 ;
        RECT 0.135 1.315 1.920 1.485 ;
        RECT 1.920 1.010 2.060 1.485 ;
        RECT 2.060 1.315 2.310 1.485 ;
        RECT 2.310 0.885 2.445 1.485 ;
        RECT 2.445 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.340 0.390 ;
        RECT 0.340 -0.085 1.940 0.085 ;
        RECT 1.940 -0.085 2.095 0.310 ;
        RECT 2.095 -0.085 2.325 0.085 ;
        RECT 2.325 -0.085 2.460 0.310 ;
        RECT 2.460 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.135 0.530 ;
      RECT 0.135 0.455 0.410 0.530 ;
      RECT 0.410 0.310 0.480 0.530 ;
      RECT 0.480 0.310 1.595 0.380 ;
      RECT 1.595 0.310 1.720 0.600 ;
      RECT 1.080 1.145 1.720 1.225 ;
      RECT 0.815 0.175 1.785 0.245 ;
      RECT 1.720 0.530 1.785 0.600 ;
      RECT 0.815 1.010 1.785 1.080 ;
      RECT 1.785 0.530 1.855 1.080 ;
      RECT 1.785 0.175 1.875 0.345 ;
      RECT 1.920 0.745 2.125 0.945 ;
      RECT 2.125 0.745 2.215 1.165 ;
      RECT 1.855 0.530 2.270 0.655 ;
      RECT 1.970 0.375 2.335 0.465 ;
      RECT 2.215 0.745 2.335 0.820 ;
      RECT 2.335 0.375 2.405 0.820 ;
  END
END NCL3W3111OF4X2

MACRO NCL4W1111OF4X1
  CLASS CORE ;
  FOREIGN NCL4W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.110 0.595 0.665 0.805 ;
        RECT 0.665 0.715 0.960 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.455 0.970 0.530 ;
        RECT 0.970 0.320 1.150 0.530 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.870 1.145 0.960 ;
        RECT 1.145 0.595 1.235 0.960 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 1.570 0.590 1.890 0.680 ;
        RECT 1.890 0.590 2.100 0.830 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 2.525 0.245 2.615 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.245 1.485 ;
        RECT 0.245 1.175 0.380 1.485 ;
        RECT 0.380 1.315 0.605 1.485 ;
        RECT 0.605 1.175 0.770 1.485 ;
        RECT 0.770 1.315 2.005 1.485 ;
        RECT 2.005 1.035 2.100 1.485 ;
        RECT 2.100 1.315 2.355 1.485 ;
        RECT 2.355 0.620 2.445 1.485 ;
        RECT 2.445 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.215 0.085 ;
        RECT 0.215 -0.085 0.380 0.255 ;
        RECT 0.380 -0.085 0.605 0.085 ;
        RECT 0.605 -0.085 0.770 0.255 ;
        RECT 0.770 -0.085 1.965 0.085 ;
        RECT 1.965 -0.085 2.060 0.255 ;
        RECT 2.060 -0.085 2.355 0.085 ;
        RECT 2.355 -0.085 2.445 0.450 ;
        RECT 2.445 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.160 0.145 0.390 ;
      RECT 0.045 1.035 0.180 1.240 ;
      RECT 0.145 0.320 0.445 0.390 ;
      RECT 0.445 0.160 0.540 0.390 ;
      RECT 0.540 0.320 0.835 0.390 ;
      RECT 0.835 0.175 0.905 0.390 ;
      RECT 1.300 0.320 1.370 0.970 ;
      RECT 1.435 0.455 1.505 0.815 ;
      RECT 1.370 0.880 1.690 0.970 ;
      RECT 1.505 0.745 1.755 0.815 ;
      RECT 1.755 0.745 1.825 0.970 ;
      RECT 0.905 0.175 1.900 0.255 ;
      RECT 0.180 1.035 1.935 1.110 ;
      RECT 1.370 0.320 2.135 0.390 ;
      RECT 1.825 0.895 2.165 0.970 ;
      RECT 1.505 0.455 2.200 0.525 ;
      RECT 2.200 0.160 2.290 0.525 ;
      RECT 2.165 0.895 2.290 1.195 ;
  END
END NCL4W1111OF4X1

MACRO NCL4W1111OF4X2
  CLASS CORE ;
  FOREIGN NCL4W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.090 0.450 0.390 0.670 ;
        RECT 0.390 0.590 0.960 0.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.545 0.435 1.170 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.735 0.940 0.805 ;
        RECT 0.940 0.735 1.080 1.085 ;
        RECT 1.080 0.590 1.170 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 1.370 0.525 1.470 0.825 ;
        RECT 1.470 0.735 1.925 0.825 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079750 ;
    PORT
      LAYER metal1 ;
        RECT 2.165 0.525 2.335 0.645 ;
        RECT 2.335 0.170 2.425 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.200 1.485 ;
        RECT 0.200 1.005 0.335 1.485 ;
        RECT 0.335 1.315 0.585 1.485 ;
        RECT 0.585 1.005 0.720 1.485 ;
        RECT 0.720 1.315 1.785 1.485 ;
        RECT 1.785 0.945 1.925 1.485 ;
        RECT 1.925 1.315 2.165 1.485 ;
        RECT 2.165 0.710 2.255 1.485 ;
        RECT 2.255 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.335 0.235 ;
        RECT 0.335 -0.085 0.585 0.085 ;
        RECT 0.585 -0.085 0.720 0.235 ;
        RECT 0.720 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.925 0.245 ;
        RECT 1.925 -0.085 2.165 0.085 ;
        RECT 2.165 -0.085 2.255 0.450 ;
        RECT 2.255 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.170 0.135 0.370 ;
      RECT 0.045 0.870 0.135 1.210 ;
      RECT 0.135 0.300 0.400 0.370 ;
      RECT 0.135 0.870 0.400 0.940 ;
      RECT 0.400 0.170 0.520 0.370 ;
      RECT 0.400 0.870 0.520 1.210 ;
      RECT 0.520 0.300 0.790 0.370 ;
      RECT 0.520 0.870 0.790 0.940 ;
      RECT 0.790 0.870 0.860 1.220 ;
      RECT 0.790 0.175 0.960 0.370 ;
      RECT 1.235 0.310 1.305 0.960 ;
      RECT 1.305 0.890 1.370 0.960 ;
      RECT 1.370 0.890 1.470 1.050 ;
      RECT 0.860 1.150 1.535 1.220 ;
      RECT 1.535 0.450 1.670 0.670 ;
      RECT 0.960 0.175 1.720 0.245 ;
      RECT 1.535 0.945 1.720 1.220 ;
      RECT 1.305 0.310 1.785 0.385 ;
      RECT 1.785 0.310 1.945 0.535 ;
      RECT 1.670 0.600 2.010 0.670 ;
      RECT 2.010 0.170 2.100 1.210 ;
  END
END NCL4W1111OF4X2

MACRO NCL4W1111OF4X4
  CLASS CORE ;
  FOREIGN NCL4W1111OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051250 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.540 0.390 0.810 ;
        RECT 0.390 0.730 0.820 0.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.540 1.150 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052250 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.875 0.915 0.965 ;
        RECT 0.915 0.785 1.215 0.965 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 1.305 0.735 1.765 0.825 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.159500 ;
    PORT
      LAYER metal1 ;
        RECT 2.120 0.540 2.315 0.905 ;
        RECT 2.315 0.540 2.580 0.810 ;
        RECT 2.580 0.540 2.595 0.910 ;
        RECT 2.595 0.370 2.670 0.910 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.220 1.485 ;
        RECT 0.220 1.240 0.355 1.485 ;
        RECT 0.355 1.315 0.615 1.485 ;
        RECT 0.615 1.240 0.820 1.485 ;
        RECT 0.820 1.315 1.815 1.485 ;
        RECT 1.815 1.095 1.935 1.485 ;
        RECT 1.935 1.315 2.305 1.485 ;
        RECT 2.305 1.160 2.510 1.485 ;
        RECT 2.510 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.220 0.085 ;
        RECT 0.220 -0.085 0.355 0.250 ;
        RECT 0.355 -0.085 0.615 0.085 ;
        RECT 0.615 -0.085 0.820 0.250 ;
        RECT 0.820 -0.085 1.895 0.085 ;
        RECT 1.895 -0.085 1.985 0.285 ;
        RECT 1.985 -0.085 2.305 0.085 ;
        RECT 2.305 -0.085 2.395 0.280 ;
        RECT 2.395 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.055 0.175 0.145 0.415 ;
      RECT 0.045 0.985 0.150 1.155 ;
      RECT 0.145 0.335 0.445 0.415 ;
      RECT 0.445 0.175 0.525 0.415 ;
      RECT 1.280 0.480 1.530 0.645 ;
      RECT 0.525 0.340 1.610 0.415 ;
      RECT 1.610 0.340 1.690 0.475 ;
      RECT 0.150 1.075 1.725 1.155 ;
      RECT 1.385 0.175 1.755 0.255 ;
      RECT 1.755 0.175 1.830 0.450 ;
      RECT 1.530 0.565 1.855 0.645 ;
      RECT 1.305 0.920 1.855 1.010 ;
      RECT 1.855 0.565 1.935 1.010 ;
      RECT 1.935 0.565 2.030 0.900 ;
      RECT 1.830 0.370 2.075 0.450 ;
      RECT 2.025 0.990 2.160 1.195 ;
      RECT 2.075 0.175 2.210 0.450 ;
      RECT 2.210 0.370 2.460 0.450 ;
      RECT 2.460 0.175 2.530 0.450 ;
      RECT 2.530 0.175 2.735 0.280 ;
      RECT 2.160 0.990 2.735 1.070 ;
      RECT 2.735 0.175 2.805 1.070 ;
  END
END NCL4W1111OF4X4

MACRO NCLAO22OF4X1
  CLASS CORE ;
  FOREIGN NCLAO22OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.595 1.700 0.665 ;
        RECT 1.700 0.595 1.715 0.810 ;
        RECT 1.715 0.535 1.955 0.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.445 1.545 0.530 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.315 0.730 0.730 0.810 ;
        RECT 0.730 0.595 1.005 0.810 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.310 0.580 0.665 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.510 0.535 2.715 0.625 ;
        RECT 2.715 0.245 2.805 0.935 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 1.035 1.485 ;
        RECT 1.035 1.290 1.175 1.485 ;
        RECT 1.175 1.315 2.160 1.485 ;
        RECT 2.160 1.000 2.395 1.485 ;
        RECT 2.395 1.315 2.510 1.485 ;
        RECT 2.510 0.690 2.645 1.485 ;
        RECT 2.645 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.115 0.295 ;
        RECT 0.115 -0.085 1.880 0.085 ;
        RECT 1.880 -0.085 2.095 0.175 ;
        RECT 2.095 -0.085 2.510 0.085 ;
        RECT 2.510 -0.085 2.645 0.470 ;
        RECT 2.645 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.930 0.115 1.225 ;
      RECT 0.180 0.175 0.250 0.945 ;
      RECT 0.250 0.875 0.400 0.945 ;
      RECT 0.400 0.875 0.490 1.090 ;
      RECT 0.115 1.155 0.555 1.225 ;
      RECT 0.555 0.875 0.625 1.225 ;
      RECT 0.250 0.175 0.645 0.245 ;
      RECT 0.645 0.175 0.715 0.380 ;
      RECT 0.625 0.875 1.070 0.945 ;
      RECT 1.070 0.730 1.140 0.945 ;
      RECT 0.875 1.010 1.205 1.090 ;
      RECT 1.205 0.875 1.275 1.090 ;
      RECT 1.140 0.730 1.580 0.810 ;
      RECT 0.715 0.310 1.610 0.380 ;
      RECT 1.610 0.310 1.680 0.470 ;
      RECT 0.780 0.175 1.745 0.245 ;
      RECT 1.745 0.175 1.815 0.335 ;
      RECT 0.690 1.155 1.885 1.225 ;
      RECT 1.680 0.400 2.020 0.470 ;
      RECT 1.275 0.875 2.020 0.945 ;
      RECT 2.020 0.400 2.095 0.945 ;
      RECT 1.510 1.010 2.095 1.090 ;
      RECT 1.815 0.265 2.160 0.335 ;
      RECT 2.095 0.535 2.290 0.670 ;
      RECT 2.160 0.400 2.355 0.470 ;
      RECT 2.160 0.155 2.395 0.335 ;
      RECT 2.355 0.400 2.445 0.935 ;
  END
END NCLAO22OF4X1

MACRO NCLAO22OF4X2
  CLASS CORE ;
  FOREIGN NCLAO22OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 3.230 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 1.225 0.590 2.330 0.675 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.455 1.925 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050750 ;
    PORT
      LAYER metal1 ;
        RECT 0.360 0.455 1.025 0.525 ;
        RECT 1.025 0.455 1.160 0.675 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050750 ;
    PORT
      LAYER metal1 ;
        RECT 0.340 0.590 0.960 0.675 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.077550 ;
    PORT
      LAYER metal1 ;
        RECT 3.095 0.230 3.185 1.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.995 1.485 ;
        RECT 0.995 1.280 1.275 1.485 ;
        RECT 1.275 1.315 2.550 1.485 ;
        RECT 2.550 1.005 2.650 1.485 ;
        RECT 2.650 1.315 2.925 1.485 ;
        RECT 2.925 0.620 3.015 1.485 ;
        RECT 3.015 1.315 3.230 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.140 0.325 ;
        RECT 0.140 -0.085 2.260 0.085 ;
        RECT 2.260 -0.085 2.485 0.255 ;
        RECT 2.485 -0.085 2.895 0.085 ;
        RECT 2.895 -0.085 3.015 0.445 ;
        RECT 3.015 -0.085 3.230 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.865 0.135 1.215 ;
      RECT 0.205 0.300 0.275 0.940 ;
      RECT 0.275 0.805 0.395 0.940 ;
      RECT 0.395 0.805 0.490 1.080 ;
      RECT 0.135 1.145 0.555 1.215 ;
      RECT 0.555 0.740 0.625 1.215 ;
      RECT 0.690 0.875 0.780 1.215 ;
      RECT 0.275 0.300 0.865 0.390 ;
      RECT 0.915 0.175 1.060 0.255 ;
      RECT 0.865 0.320 1.095 0.390 ;
      RECT 1.095 0.310 1.275 0.390 ;
      RECT 1.060 0.175 1.310 0.245 ;
      RECT 1.310 0.175 1.480 0.255 ;
      RECT 1.275 0.320 1.515 0.390 ;
      RECT 0.625 0.740 1.670 0.810 ;
      RECT 1.515 0.310 1.990 0.390 ;
      RECT 1.990 0.310 2.060 0.525 ;
      RECT 1.480 0.175 2.125 0.245 ;
      RECT 2.125 0.175 2.195 0.390 ;
      RECT 0.780 1.145 2.290 1.215 ;
      RECT 1.685 1.010 2.355 1.080 ;
      RECT 2.060 0.455 2.410 0.525 ;
      RECT 0.845 0.875 2.410 0.945 ;
      RECT 2.410 0.455 2.480 0.945 ;
      RECT 2.355 1.010 2.485 1.250 ;
      RECT 2.195 0.320 2.550 0.390 ;
      RECT 2.550 0.230 2.650 0.390 ;
      RECT 2.480 0.455 2.675 0.590 ;
      RECT 2.545 0.655 2.740 0.940 ;
      RECT 2.740 0.320 2.830 0.940 ;
  END
END NCLAO22OF4X2

MACRO NCLAO22OF4X4
  CLASS CORE ;
  FOREIGN NCLAO22OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 3.230 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050750 ;
    PORT
      LAYER metal1 ;
        RECT 0.155 0.460 0.380 0.675 ;
        RECT 0.380 0.595 0.770 0.675 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.470 0.445 0.960 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.030 0.730 1.135 0.965 ;
        RECT 1.135 0.730 1.725 0.815 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.450 1.340 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.206900 ;
    PORT
      LAYER metal1 ;
        RECT 2.720 0.755 2.800 1.225 ;
        RECT 2.555 0.290 3.080 0.370 ;
        RECT 3.080 0.165 3.095 0.370 ;
        RECT 2.800 0.755 3.095 0.835 ;
        RECT 3.095 0.165 3.115 0.835 ;
        RECT 3.115 0.165 3.185 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.515 1.485 ;
        RECT 0.515 1.055 0.745 1.485 ;
        RECT 0.745 1.315 2.370 1.485 ;
        RECT 2.370 1.050 2.460 1.485 ;
        RECT 2.460 1.315 2.890 1.485 ;
        RECT 2.890 0.915 3.025 1.485 ;
        RECT 3.025 1.315 3.230 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.285 0.260 ;
        RECT 0.285 -0.085 1.810 0.085 ;
        RECT 1.810 -0.085 1.945 0.165 ;
        RECT 1.945 -0.085 2.195 0.085 ;
        RECT 2.195 -0.085 2.285 0.370 ;
        RECT 2.285 -0.085 2.760 0.085 ;
        RECT 2.760 -0.085 2.990 0.200 ;
        RECT 2.990 -0.085 3.230 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.755 0.125 1.090 ;
      RECT 0.470 0.220 0.610 0.380 ;
      RECT 0.125 0.755 0.860 0.835 ;
      RECT 0.205 0.905 0.860 0.985 ;
      RECT 0.860 0.595 0.940 0.835 ;
      RECT 0.860 0.905 0.940 1.205 ;
      RECT 0.610 0.310 1.430 0.380 ;
      RECT 1.430 0.310 1.530 0.505 ;
      RECT 0.940 1.055 1.580 1.205 ;
      RECT 0.700 0.175 1.640 0.245 ;
      RECT 1.280 0.905 1.645 0.985 ;
      RECT 1.640 0.175 1.720 0.335 ;
      RECT 1.645 0.905 1.725 1.225 ;
      RECT 0.940 0.595 1.800 0.665 ;
      RECT 1.800 0.595 1.870 1.090 ;
      RECT 1.530 0.425 1.935 0.505 ;
      RECT 1.935 0.425 2.015 0.950 ;
      RECT 1.720 0.255 2.105 0.335 ;
      RECT 1.870 1.015 2.160 1.090 ;
      RECT 2.015 0.755 2.225 0.950 ;
      RECT 1.725 1.155 2.225 1.225 ;
      RECT 2.225 0.755 2.305 1.225 ;
      RECT 2.105 0.460 2.375 0.665 ;
      RECT 2.305 0.755 2.460 0.960 ;
      RECT 2.375 0.290 2.465 0.665 ;
      RECT 2.465 0.465 2.550 0.665 ;
      RECT 2.550 0.465 2.630 1.185 ;
      RECT 2.720 0.460 2.940 0.665 ;
  END
END NCLAO22OF4X4

MACRO NCLOA22OF4X1
  CLASS CORE ;
  FOREIGN NCLOA22OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.735 1.510 0.805 ;
        RECT 1.510 0.735 1.720 0.945 ;
        RECT 1.720 0.735 2.355 0.805 ;
        RECT 2.355 0.610 2.490 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.595 1.990 0.670 ;
        RECT 1.990 0.455 2.290 0.670 ;
        RECT 2.290 0.455 2.490 0.545 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.870 1.445 0.955 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.455 1.910 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.041800 ;
    PORT
      LAYER metal1 ;
        RECT 2.715 0.175 2.805 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.240 1.485 ;
        RECT 0.240 0.930 0.330 1.485 ;
        RECT 0.330 1.315 2.355 1.485 ;
        RECT 2.355 1.035 2.650 1.485 ;
        RECT 2.650 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.330 0.255 ;
        RECT 0.330 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.225 0.110 ;
        RECT 2.225 -0.085 2.520 0.085 ;
        RECT 2.520 -0.085 2.610 0.255 ;
        RECT 2.610 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.135 1.190 ;
      RECT 0.135 0.660 0.345 0.865 ;
      RECT 0.200 0.320 0.425 0.595 ;
      RECT 0.425 0.320 0.495 1.090 ;
      RECT 0.495 1.020 1.090 1.090 ;
      RECT 0.395 0.175 1.470 0.255 ;
      RECT 0.560 1.155 1.515 1.225 ;
      RECT 0.495 0.320 1.535 0.390 ;
      RECT 1.535 0.230 1.660 0.390 ;
      RECT 1.535 1.010 2.225 1.090 ;
      RECT 1.725 0.175 2.450 0.255 ;
      RECT 1.660 0.320 2.560 0.390 ;
      RECT 1.925 0.870 2.560 0.945 ;
      RECT 2.560 0.320 2.650 0.945 ;
  END
END NCLOA22OF4X1

MACRO NCLOA22OF4X2
  CLASS CORE ;
  FOREIGN NCLOA22OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 0.655 0.515 0.755 1.040 ;
        RECT 0.755 0.515 0.805 0.945 ;
        RECT 0.805 0.875 2.325 0.945 ;
        RECT 2.325 0.515 2.480 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050500 ;
    PORT
      LAYER metal1 ;
        RECT 0.915 0.730 2.260 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.455 1.720 0.530 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.595 1.860 0.665 ;
        RECT 1.860 0.455 2.160 0.665 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079750 ;
    PORT
      LAYER metal1 ;
        RECT 2.715 0.150 2.805 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.285 1.485 ;
        RECT 0.285 0.920 0.495 1.485 ;
        RECT 0.495 1.315 2.430 1.485 ;
        RECT 2.430 1.145 2.610 1.485 ;
        RECT 2.610 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.235 0.085 ;
        RECT 0.235 -0.085 0.330 0.245 ;
        RECT 0.330 -0.085 2.005 0.085 ;
        RECT 2.005 -0.085 2.235 0.120 ;
        RECT 2.235 -0.085 2.515 0.085 ;
        RECT 2.515 -0.085 2.610 0.200 ;
        RECT 2.610 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.115 1.185 ;
      RECT 0.115 0.650 0.135 1.185 ;
      RECT 0.180 0.310 0.285 0.585 ;
      RECT 0.135 0.650 0.590 0.855 ;
      RECT 0.395 0.175 1.485 0.245 ;
      RECT 0.585 1.145 1.485 1.225 ;
      RECT 0.285 0.310 1.550 0.390 ;
      RECT 1.550 0.220 1.670 0.390 ;
      RECT 1.550 1.145 2.235 1.225 ;
      RECT 1.735 0.185 2.450 0.255 ;
      RECT 1.670 0.320 2.570 0.390 ;
      RECT 0.970 1.010 2.570 1.080 ;
      RECT 2.570 0.320 2.650 1.080 ;
  END
END NCLOA22OF4X2

MACRO NCLOA22OF4X4
  CLASS CORE ;
  FOREIGN NCLOA22OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 3.230 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.590 2.035 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.200 0.665 0.280 1.090 ;
        RECT 0.280 1.015 1.025 1.090 ;
        RECT 1.025 0.870 1.105 1.090 ;
        RECT 1.105 0.870 1.670 0.940 ;
        RECT 1.670 0.755 1.805 0.940 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.480 0.730 1.580 0.805 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.870 0.960 0.950 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 2.895 0.245 2.990 1.160 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 1.880 1.485 ;
        RECT 1.880 1.290 2.160 1.485 ;
        RECT 2.160 1.315 2.715 1.485 ;
        RECT 2.715 0.945 2.805 1.485 ;
        RECT 2.805 1.315 3.095 1.485 ;
        RECT 3.095 0.805 3.185 1.485 ;
        RECT 3.185 1.315 3.230 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.225 0.085 ;
        RECT 0.225 -0.085 0.360 0.185 ;
        RECT 0.360 -0.085 2.380 0.085 ;
        RECT 2.380 -0.085 2.470 0.310 ;
        RECT 2.470 -0.085 2.715 0.085 ;
        RECT 2.715 -0.085 2.805 0.455 ;
        RECT 2.805 -0.085 3.095 0.085 ;
        RECT 3.095 -0.085 3.185 0.445 ;
        RECT 3.185 -0.085 3.230 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.445 0.125 1.230 ;
      RECT 0.045 0.175 0.135 0.355 ;
      RECT 0.135 0.275 0.450 0.355 ;
      RECT 0.450 0.175 0.535 0.355 ;
      RECT 0.125 0.445 0.625 0.525 ;
      RECT 0.625 0.345 0.790 0.525 ;
      RECT 0.535 0.175 0.870 0.255 ;
      RECT 0.870 0.175 0.950 0.345 ;
      RECT 0.790 0.435 1.025 0.525 ;
      RECT 1.025 0.175 1.105 0.525 ;
      RECT 0.420 1.155 1.270 1.225 ;
      RECT 1.105 0.455 2.100 0.525 ;
      RECT 1.170 1.005 2.100 1.075 ;
      RECT 1.170 0.310 2.175 0.390 ;
      RECT 2.100 0.455 2.180 1.075 ;
      RECT 1.105 0.175 2.245 0.245 ;
      RECT 2.245 0.175 2.315 0.835 ;
      RECT 1.270 1.145 2.385 1.225 ;
      RECT 2.315 0.630 2.445 0.835 ;
      RECT 2.395 0.400 2.535 0.540 ;
      RECT 2.535 0.400 2.625 1.220 ;
  END
END NCLOA22OF4X4

MACRO NCLP1W1111OF4X1
  CLASS CORE ;
  FOREIGN NCLP1W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.535 0.455 0.795 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.505 0.730 0.795 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.455 0.470 0.530 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.595 0.390 0.900 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 1.010 0.230 1.095 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.970 0.135 1.485 ;
        RECT 0.135 1.315 0.415 1.485 ;
        RECT 0.415 1.145 0.550 1.485 ;
        RECT 0.550 1.315 0.800 1.485 ;
        RECT 0.800 1.145 0.945 1.485 ;
        RECT 0.945 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.725 0.085 ;
        RECT 0.725 -0.085 0.945 0.255 ;
        RECT 0.945 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.115 0.480 ;
      RECT 0.115 0.150 0.135 0.390 ;
      RECT 0.210 1.010 0.350 1.250 ;
      RECT 0.350 1.010 0.625 1.080 ;
      RECT 0.625 1.010 0.715 1.250 ;
      RECT 0.135 0.320 0.870 0.390 ;
      RECT 0.715 1.010 0.870 1.080 ;
      RECT 0.870 0.320 0.945 1.080 ;
  END
END NCLP1W1111OF4X1

MACRO NCLP1W1111OF4X2
  CLASS CORE ;
  FOREIGN NCLP1W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.790 0.245 0.890 0.620 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.410 0.245 0.700 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.800 0.770 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.205 0.245 0.320 0.735 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.005 0.170 1.095 1.230 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.050 1.485 ;
        RECT 0.050 1.170 0.140 1.485 ;
        RECT 0.140 1.315 0.410 1.485 ;
        RECT 0.410 1.185 0.545 1.485 ;
        RECT 0.545 1.315 0.800 1.485 ;
        RECT 0.800 1.185 0.940 1.485 ;
        RECT 0.940 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.800 0.085 ;
        RECT 0.800 -0.085 0.940 0.180 ;
        RECT 0.940 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.220 0.115 1.105 ;
      RECT 0.115 1.035 0.210 1.105 ;
      RECT 0.210 1.035 0.345 1.230 ;
      RECT 0.345 1.035 0.610 1.105 ;
      RECT 0.610 1.035 0.735 1.230 ;
      RECT 0.735 1.035 0.850 1.105 ;
      RECT 0.850 0.690 0.940 1.105 ;
  END
END NCLP1W1111OF4X2

MACRO NCLP1W1111OF4X4
  CLASS CORE ;
  FOREIGN NCLP1W1111OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.330 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.735 0.785 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 0.600 0.385 0.710 0.660 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 0.315 0.385 0.510 0.595 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.665 0.390 0.945 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.102200 ;
    PORT
      LAYER metal1 ;
        RECT 1.010 0.175 1.100 1.235 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.060 1.485 ;
        RECT 0.060 1.030 0.140 1.485 ;
        RECT 0.140 1.315 0.455 1.485 ;
        RECT 0.455 1.170 0.535 1.485 ;
        RECT 0.535 1.315 0.840 1.485 ;
        RECT 0.840 1.170 0.920 1.485 ;
        RECT 0.920 1.315 1.195 1.485 ;
        RECT 1.195 0.830 1.285 1.485 ;
        RECT 1.285 1.315 1.330 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.800 0.085 ;
        RECT 0.800 -0.085 0.935 0.185 ;
        RECT 0.935 -0.085 1.195 0.085 ;
        RECT 1.195 -0.085 1.285 0.430 ;
        RECT 1.285 -0.085 1.330 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.180 0.430 ;
      RECT 0.230 1.010 0.365 1.225 ;
      RECT 0.365 1.010 0.615 1.090 ;
      RECT 0.180 0.175 0.630 0.255 ;
      RECT 0.630 0.175 0.710 0.320 ;
      RECT 0.615 1.010 0.750 1.225 ;
      RECT 0.710 0.250 0.865 0.320 ;
      RECT 0.750 1.010 0.865 1.090 ;
      RECT 0.865 0.250 0.945 1.090 ;
  END
END NCLP1W1111OF4X4

MACRO NCLP1W111OF3X1
  CLASS CORE ;
  FOREIGN NCLP1W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.605 0.600 0.880 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.315 0.440 0.540 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.640 0.360 0.880 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 0.815 0.245 0.905 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.250 1.485 ;
        RECT 0.250 1.080 0.360 1.485 ;
        RECT 0.360 1.315 0.640 1.485 ;
        RECT 0.640 1.085 0.745 1.485 ;
        RECT 0.745 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.640 0.085 ;
        RECT 0.640 -0.085 0.745 0.370 ;
        RECT 0.745 -0.085 0.950 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.115 0.450 ;
      RECT 0.045 0.945 0.175 1.225 ;
      RECT 0.175 0.945 0.440 1.015 ;
      RECT 0.115 0.175 0.505 0.250 ;
      RECT 0.440 0.945 0.540 1.225 ;
      RECT 0.505 0.175 0.575 0.505 ;
      RECT 0.575 0.435 0.670 0.505 ;
      RECT 0.540 0.945 0.670 1.020 ;
      RECT 0.670 0.435 0.745 1.020 ;
  END
END NCLP1W111OF3X1

MACRO NCLP1W111OF3X2
  CLASS CORE ;
  FOREIGN NCLP1W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020500 ;
    PORT
      LAYER metal1 ;
        RECT 0.495 0.390 0.595 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020500 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.390 0.405 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020500 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.595 0.390 0.805 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 0.820 0.175 0.905 1.110 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.215 1.485 ;
        RECT 0.215 1.065 0.350 1.485 ;
        RECT 0.350 1.315 0.605 1.485 ;
        RECT 0.605 1.065 0.740 1.485 ;
        RECT 0.740 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.585 0.085 ;
        RECT 0.585 -0.085 0.720 0.160 ;
        RECT 0.720 -0.085 0.950 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.895 0.125 1.065 ;
      RECT 0.125 0.895 0.440 0.975 ;
      RECT 0.045 0.175 0.495 0.310 ;
      RECT 0.440 0.895 0.520 1.065 ;
      RECT 0.495 0.230 0.675 0.310 ;
      RECT 0.520 0.895 0.675 0.975 ;
      RECT 0.675 0.230 0.755 0.975 ;
  END
END NCLP1W111OF3X2

MACRO NCLP1W111OF3X4
  CLASS CORE ;
  FOREIGN NCLP1W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.140 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.435 0.625 0.595 0.900 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.400 0.405 0.535 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.020750 ;
    PORT
      LAYER metal1 ;
        RECT 0.145 0.625 0.345 0.875 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 0.820 0.175 0.910 1.070 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.210 1.485 ;
        RECT 0.210 1.160 0.345 1.485 ;
        RECT 0.345 1.315 0.605 1.485 ;
        RECT 0.605 1.160 0.745 1.485 ;
        RECT 0.745 1.315 1.005 1.485 ;
        RECT 1.005 0.845 1.095 1.485 ;
        RECT 1.095 1.315 1.140 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.640 0.085 ;
        RECT 0.640 -0.085 0.730 0.365 ;
        RECT 0.730 -0.085 1.005 0.085 ;
        RECT 1.005 -0.085 1.095 0.365 ;
        RECT 1.095 -0.085 1.140 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.990 0.125 1.160 ;
      RECT 0.125 0.990 0.435 1.070 ;
      RECT 0.045 0.175 0.470 0.310 ;
      RECT 0.435 0.990 0.515 1.160 ;
      RECT 0.470 0.175 0.550 0.535 ;
      RECT 0.550 0.455 0.665 0.535 ;
      RECT 0.515 0.990 0.665 1.070 ;
      RECT 0.665 0.455 0.745 1.070 ;
  END
END NCLP1W111OF3X4

MACRO NCLP1W11OF2X1
  CLASS CORE ;
  FOREIGN NCLP1W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.595 0.395 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.395 0.410 0.530 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.170 0.715 1.215 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.940 0.135 1.485 ;
        RECT 0.135 1.315 0.420 1.485 ;
        RECT 0.420 1.110 0.560 1.485 ;
        RECT 0.560 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.560 0.195 ;
        RECT 0.560 -0.085 0.760 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.170 0.180 0.330 ;
      RECT 0.220 0.970 0.355 1.180 ;
      RECT 0.180 0.260 0.475 0.330 ;
      RECT 0.355 0.970 0.475 1.040 ;
      RECT 0.475 0.260 0.560 1.040 ;
  END
END NCLP1W11OF2X1

MACRO NCLP1W11OF2X2
  CLASS CORE ;
  FOREIGN NCLP1W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.760 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.160 0.730 0.400 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.425 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078100 ;
    PORT
      LAYER metal1 ;
        RECT 0.625 0.150 0.715 1.230 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.005 0.130 1.485 ;
        RECT 0.130 1.315 0.420 1.485 ;
        RECT 0.420 1.145 0.560 1.485 ;
        RECT 0.560 1.315 0.760 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.560 0.160 ;
        RECT 0.560 -0.085 0.760 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.190 0.295 ;
      RECT 0.220 1.010 0.355 1.250 ;
      RECT 0.190 0.225 0.490 0.295 ;
      RECT 0.355 1.010 0.490 1.080 ;
      RECT 0.490 0.225 0.560 1.080 ;
  END
END NCLP1W11OF2X2

MACRO NCLP1W11OF2X4
  CLASS CORE ;
  FOREIGN NCLP1W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.950 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.180 0.595 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.019750 ;
    PORT
      LAYER metal1 ;
        RECT 0.175 0.665 0.405 0.805 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.102950 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.175 0.720 1.110 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.895 0.135 1.485 ;
        RECT 0.135 1.315 0.410 1.485 ;
        RECT 0.410 1.065 0.545 1.485 ;
        RECT 0.545 1.315 0.810 1.485 ;
        RECT 0.810 0.705 0.900 1.485 ;
        RECT 0.900 1.315 0.950 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.440 0.085 ;
        RECT 0.440 -0.085 0.540 0.235 ;
        RECT 0.540 -0.085 0.810 0.085 ;
        RECT 0.810 -0.085 0.900 0.375 ;
        RECT 0.900 -0.085 0.950 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.270 0.310 ;
      RECT 0.225 0.895 0.320 1.170 ;
      RECT 0.270 0.175 0.350 0.405 ;
      RECT 0.350 0.325 0.485 0.405 ;
      RECT 0.320 0.895 0.485 0.975 ;
      RECT 0.485 0.325 0.565 0.975 ;
  END
END NCLP1W11OF2X4

MACRO NCLP2W11OF2X1
  CLASS CORE ;
  FOREIGN NCLP2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.710 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.041750 ;
    PORT
      LAYER metal1 ;
        RECT 0.170 0.805 0.710 1.015 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.041750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.510 0.960 0.715 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 1.360 0.385 1.575 0.685 ;
        RECT 1.575 0.155 1.665 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.065 0.125 1.485 ;
        RECT 0.125 1.315 0.395 1.485 ;
        RECT 0.395 1.240 0.540 1.485 ;
        RECT 0.540 1.315 1.380 1.485 ;
        RECT 1.380 0.820 1.470 1.485 ;
        RECT 1.470 1.315 1.710 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.050 0.085 ;
        RECT 0.050 -0.085 0.140 0.400 ;
        RECT 0.140 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.540 0.280 ;
        RECT 0.540 -0.085 1.360 0.085 ;
        RECT 1.360 -0.085 1.470 0.310 ;
        RECT 1.470 -0.085 1.710 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.255 0.310 0.415 ;
      RECT 0.205 1.105 0.605 1.175 ;
      RECT 0.310 0.345 0.640 0.415 ;
      RECT 0.605 1.105 0.675 1.225 ;
      RECT 0.640 0.175 0.710 0.415 ;
      RECT 0.780 0.310 0.940 0.445 ;
      RECT 0.780 0.780 0.940 1.070 ;
      RECT 0.710 0.175 1.005 0.245 ;
      RECT 0.675 1.155 1.005 1.225 ;
      RECT 0.940 0.375 1.050 0.445 ;
      RECT 0.940 0.780 1.050 0.955 ;
      RECT 1.005 0.175 1.140 0.310 ;
      RECT 1.050 0.375 1.140 0.955 ;
      RECT 1.005 1.020 1.140 1.225 ;
      RECT 1.205 0.155 1.295 1.225 ;
  END
END NCLP2W11OF2X1

MACRO NCLP2W11OF2X2
  CLASS CORE ;
  FOREIGN NCLP2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.730 0.820 0.820 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.042000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.575 0.995 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.520 0.440 1.765 0.740 ;
        RECT 1.765 0.245 1.855 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.055 1.485 ;
        RECT 0.055 0.885 0.150 1.485 ;
        RECT 0.150 1.315 0.400 1.485 ;
        RECT 0.400 1.040 0.685 1.485 ;
        RECT 0.685 1.315 1.520 1.485 ;
        RECT 1.520 0.885 1.660 1.485 ;
        RECT 1.660 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.070 0.085 ;
        RECT 0.070 -0.085 0.180 0.430 ;
        RECT 0.180 -0.085 0.425 0.085 ;
        RECT 0.425 -0.085 0.595 0.370 ;
        RECT 0.595 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.660 0.365 ;
        RECT 1.660 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.245 0.300 0.360 0.510 ;
      RECT 0.360 0.440 0.660 0.510 ;
      RECT 0.660 0.175 0.735 0.510 ;
      RECT 0.215 0.885 0.750 0.975 ;
      RECT 0.750 0.885 0.820 1.225 ;
      RECT 0.805 0.335 1.060 0.510 ;
      RECT 0.885 0.730 1.060 1.090 ;
      RECT 1.060 0.335 1.100 1.090 ;
      RECT 1.100 0.335 1.130 0.855 ;
      RECT 0.820 1.155 1.165 1.225 ;
      RECT 0.735 0.175 1.195 0.245 ;
      RECT 1.195 0.175 1.300 0.430 ;
      RECT 1.130 0.555 1.300 0.855 ;
      RECT 1.165 0.920 1.300 1.225 ;
      RECT 1.365 0.245 1.455 1.155 ;
  END
END NCLP2W11OF2X2

MACRO NCLP2W11OF2X4
  CLASS CORE ;
  FOREIGN NCLP2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.735 0.370 0.825 ;
        RECT 0.370 0.735 0.590 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.043000 ;
    PORT
      LAYER metal1 ;
        RECT 0.330 0.455 0.805 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 1.565 0.175 1.660 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.970 0.125 1.485 ;
        RECT 0.125 1.315 0.395 1.485 ;
        RECT 0.395 1.160 0.535 1.485 ;
        RECT 0.535 1.315 1.385 1.485 ;
        RECT 1.385 0.745 1.475 1.485 ;
        RECT 1.475 1.315 1.765 1.485 ;
        RECT 1.765 0.675 1.855 1.485 ;
        RECT 1.855 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.305 ;
        RECT 0.135 -0.085 0.395 0.085 ;
        RECT 0.395 -0.085 0.530 0.195 ;
        RECT 0.530 -0.085 1.385 0.085 ;
        RECT 1.385 -0.085 1.475 0.455 ;
        RECT 1.475 -0.085 1.765 0.085 ;
        RECT 1.765 -0.085 1.855 0.445 ;
        RECT 1.855 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.195 0.305 0.365 ;
      RECT 0.205 1.010 0.305 1.250 ;
      RECT 0.305 0.285 0.620 0.365 ;
      RECT 0.305 1.010 0.625 1.090 ;
      RECT 0.620 0.175 0.700 0.365 ;
      RECT 0.625 1.010 0.705 1.225 ;
      RECT 0.790 0.310 0.870 0.390 ;
      RECT 0.795 0.755 0.870 1.055 ;
      RECT 0.870 0.310 0.950 1.055 ;
      RECT 0.700 0.175 1.035 0.245 ;
      RECT 0.705 1.145 1.040 1.225 ;
      RECT 1.035 0.175 1.115 0.335 ;
      RECT 0.950 0.440 1.125 0.575 ;
      RECT 1.030 0.665 1.205 0.870 ;
      RECT 1.040 0.950 1.245 1.225 ;
      RECT 1.205 0.315 1.295 0.870 ;
  END
END NCLP2W11OF2X4

MACRO NCLP2W211OF3X1
  CLASS CORE ;
  FOREIGN NCLP2W211OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 1.295 0.595 1.725 0.685 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.285 0.455 0.460 0.570 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.120 0.660 0.700 0.875 ;
        RECT 0.700 0.660 1.020 0.750 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.105 0.385 2.220 0.950 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.965 0.125 1.485 ;
        RECT 0.125 1.315 0.420 1.485 ;
        RECT 0.420 1.150 0.555 1.485 ;
        RECT 0.555 1.315 1.395 1.485 ;
        RECT 1.395 1.135 1.535 1.485 ;
        RECT 1.535 1.315 1.935 1.485 ;
        RECT 1.935 0.675 2.015 1.485 ;
        RECT 2.015 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.415 ;
        RECT 0.135 -0.085 0.450 0.085 ;
        RECT 0.450 -0.085 0.585 0.240 ;
        RECT 0.585 -0.085 1.935 0.085 ;
        RECT 1.935 -0.085 2.015 0.490 ;
        RECT 2.015 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.210 0.965 0.315 1.225 ;
      RECT 0.225 0.175 0.360 0.390 ;
      RECT 0.315 0.965 0.645 1.060 ;
      RECT 0.645 0.965 0.725 1.225 ;
      RECT 0.815 0.840 0.970 1.045 ;
      RECT 0.360 0.310 1.125 0.390 ;
      RECT 0.725 1.135 1.125 1.225 ;
      RECT 0.815 0.175 1.205 0.245 ;
      RECT 1.125 0.460 1.205 0.865 ;
      RECT 0.970 0.955 1.215 1.045 ;
      RECT 1.215 0.955 1.305 1.225 ;
      RECT 1.205 0.175 1.340 0.380 ;
      RECT 1.430 0.175 1.725 0.380 ;
      RECT 1.305 0.955 1.725 1.045 ;
      RECT 1.205 0.460 1.845 0.530 ;
      RECT 1.205 0.775 1.845 0.865 ;
  END
END NCLP2W211OF3X1

MACRO NCLP2W211OF3X2
  CLASS CORE ;
  FOREIGN NCLP2W211OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.595 1.405 0.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.485 0.890 0.735 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.645 0.340 0.945 ;
        RECT 0.340 0.825 0.855 0.945 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078100 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.460 1.955 0.555 ;
        RECT 1.955 0.245 2.045 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.065 0.125 1.485 ;
        RECT 0.125 1.315 0.405 1.485 ;
        RECT 0.405 1.225 0.545 1.485 ;
        RECT 0.545 1.315 1.545 1.485 ;
        RECT 1.545 1.035 1.635 1.485 ;
        RECT 1.635 1.315 1.770 1.485 ;
        RECT 1.770 0.645 1.860 1.485 ;
        RECT 1.860 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.415 ;
        RECT 0.125 -0.085 0.405 0.085 ;
        RECT 0.405 -0.085 0.565 0.240 ;
        RECT 0.565 -0.085 1.770 0.085 ;
        RECT 1.770 -0.085 1.860 0.310 ;
        RECT 1.860 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.205 0.175 0.340 0.395 ;
      RECT 0.210 1.045 0.620 1.135 ;
      RECT 0.620 1.045 0.700 1.225 ;
      RECT 0.790 1.010 0.960 1.090 ;
      RECT 0.960 0.460 1.040 1.090 ;
      RECT 0.340 0.320 1.095 0.395 ;
      RECT 0.700 1.155 1.095 1.225 ;
      RECT 0.790 0.175 1.160 0.255 ;
      RECT 1.040 1.015 1.180 1.090 ;
      RECT 1.160 0.175 1.295 0.385 ;
      RECT 1.040 0.460 1.385 0.530 ;
      RECT 1.180 1.015 1.455 1.230 ;
      RECT 1.385 0.180 1.525 0.530 ;
      RECT 1.130 0.875 1.590 0.950 ;
      RECT 1.590 0.245 1.680 0.950 ;
  END
END NCLP2W211OF3X2

MACRO NCLP2W211OF3X4
  CLASS CORE ;
  FOREIGN NCLP2W211OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022750 ;
    PORT
      LAYER metal1 ;
        RECT 1.385 0.900 1.520 1.225 ;
        RECT 1.520 1.005 1.720 1.225 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.525 0.890 0.750 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.175 0.665 0.350 0.945 ;
        RECT 0.350 0.840 0.980 0.945 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.102950 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.245 2.055 1.060 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.125 1.485 ;
        RECT 0.125 1.315 0.400 1.485 ;
        RECT 0.400 1.210 0.535 1.485 ;
        RECT 0.535 1.315 1.370 1.485 ;
        RECT 1.370 1.290 1.645 1.485 ;
        RECT 1.645 1.315 1.785 1.485 ;
        RECT 1.785 0.640 1.870 1.485 ;
        RECT 1.870 1.315 2.145 1.485 ;
        RECT 2.145 0.700 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.135 0.435 ;
        RECT 0.135 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.565 0.260 ;
        RECT 0.565 -0.085 1.770 0.085 ;
        RECT 1.770 -0.085 1.870 0.305 ;
        RECT 1.870 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.445 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.225 0.160 0.310 0.435 ;
      RECT 0.205 1.035 0.625 1.120 ;
      RECT 0.625 1.035 0.705 1.225 ;
      RECT 0.310 0.350 1.080 0.435 ;
      RECT 0.705 1.155 1.085 1.225 ;
      RECT 0.790 0.175 1.155 0.260 ;
      RECT 0.795 1.010 1.160 1.090 ;
      RECT 1.160 1.010 1.190 1.225 ;
      RECT 1.155 0.175 1.235 0.480 ;
      RECT 1.190 0.730 1.295 1.225 ;
      RECT 1.050 0.560 1.300 0.640 ;
      RECT 1.300 0.175 1.370 0.640 ;
      RECT 1.295 0.730 1.435 0.810 ;
      RECT 1.435 0.345 1.515 0.810 ;
      RECT 1.370 0.175 1.590 0.255 ;
      RECT 1.590 0.175 1.680 0.915 ;
  END
END NCLP2W211OF3X4

MACRO NCLP3W111OF3X1
  CLASS CORE ;
  FOREIGN NCLP3W111OF3X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.590 0.595 0.700 0.875 ;
        RECT 0.700 0.595 1.320 0.665 ;
        RECT 1.320 0.445 1.570 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048000 ;
    PORT
      LAYER metal1 ;
        RECT 0.935 0.730 1.150 0.945 ;
        RECT 1.150 0.855 1.265 0.945 ;
        RECT 1.265 0.730 1.530 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.445 1.255 0.530 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.042350 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.150 1.855 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.200 1.485 ;
        RECT 0.200 0.970 0.325 1.485 ;
        RECT 0.325 1.315 1.520 1.485 ;
        RECT 1.520 1.145 1.705 1.485 ;
        RECT 1.705 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.235 0.085 ;
        RECT 0.235 -0.085 0.345 0.330 ;
        RECT 0.345 -0.085 1.560 0.085 ;
        RECT 1.560 -0.085 1.705 0.245 ;
        RECT 1.705 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.275 0.135 0.465 ;
      RECT 0.045 0.835 0.135 1.250 ;
      RECT 0.115 0.530 0.215 0.770 ;
      RECT 0.135 0.395 0.280 0.465 ;
      RECT 0.135 0.835 0.390 0.905 ;
      RECT 0.280 0.395 0.440 0.635 ;
      RECT 0.215 0.700 0.455 0.770 ;
      RECT 0.425 0.175 0.515 0.330 ;
      RECT 0.455 0.700 0.525 1.080 ;
      RECT 0.525 1.010 0.750 1.080 ;
      RECT 0.750 0.920 0.840 1.080 ;
      RECT 0.515 0.175 0.920 0.245 ;
      RECT 0.390 1.145 0.945 1.225 ;
      RECT 0.580 0.310 0.985 0.380 ;
      RECT 0.840 1.010 1.010 1.080 ;
      RECT 1.010 1.010 1.125 1.250 ;
      RECT 0.985 0.220 1.495 0.380 ;
      RECT 1.495 0.310 1.635 0.380 ;
      RECT 1.125 1.010 1.635 1.080 ;
      RECT 1.635 0.310 1.705 1.080 ;
  END
END NCLP3W111OF3X1

MACRO NCLP3W111OF3X2
  CLASS CORE ;
  FOREIGN NCLP3W111OF3X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 1.900 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.730 1.405 0.805 ;
        RECT 1.405 0.505 1.570 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.870 1.540 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.044000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.575 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.150 1.855 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.190 1.485 ;
        RECT 0.190 1.145 0.335 1.485 ;
        RECT 0.335 1.315 1.520 1.485 ;
        RECT 1.520 1.165 1.705 1.485 ;
        RECT 1.705 1.315 1.900 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.360 0.340 ;
        RECT 0.360 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.705 0.260 ;
        RECT 1.705 -0.085 1.900 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.290 0.125 1.145 ;
      RECT 0.125 0.290 0.135 0.650 ;
      RECT 0.190 0.715 0.280 1.080 ;
      RECT 0.135 0.445 0.475 0.650 ;
      RECT 0.425 0.185 0.525 0.340 ;
      RECT 0.590 0.325 0.765 0.485 ;
      RECT 0.525 0.185 0.830 0.255 ;
      RECT 0.830 0.185 0.925 0.340 ;
      RECT 0.400 1.145 0.945 1.225 ;
      RECT 0.765 0.415 0.990 0.485 ;
      RECT 0.280 1.010 1.010 1.080 ;
      RECT 1.010 1.010 1.130 1.250 ;
      RECT 0.990 0.325 1.150 0.485 ;
      RECT 1.150 0.325 1.635 0.395 ;
      RECT 1.130 1.010 1.635 1.100 ;
      RECT 1.635 0.325 1.705 1.100 ;
  END
END NCLP3W111OF3X2

MACRO NCLP3W111OF3X4
  CLASS CORE ;
  FOREIGN NCLP3W111OF3X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.540 0.730 1.465 0.805 ;
        RECT 1.465 0.465 1.555 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.870 0.870 1.465 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046000 ;
    PORT
      LAYER metal1 ;
        RECT 0.745 0.585 1.340 0.665 ;
    END
  END C
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.107300 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.170 1.860 1.235 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.220 1.485 ;
        RECT 0.220 0.960 0.300 1.485 ;
        RECT 0.300 1.315 1.520 1.485 ;
        RECT 1.520 1.205 1.680 1.485 ;
        RECT 1.680 1.315 1.955 1.485 ;
        RECT 1.955 0.890 2.045 1.485 ;
        RECT 2.045 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.220 0.085 ;
        RECT 0.220 -0.085 0.305 0.355 ;
        RECT 0.305 -0.085 1.520 0.085 ;
        RECT 1.520 -0.085 1.660 0.205 ;
        RECT 1.660 -0.085 1.955 0.085 ;
        RECT 1.955 -0.085 2.045 0.355 ;
        RECT 2.045 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.295 0.130 0.530 ;
      RECT 0.045 0.740 0.130 1.235 ;
      RECT 0.130 0.740 0.335 0.875 ;
      RECT 0.135 0.595 0.400 0.675 ;
      RECT 0.130 0.445 0.435 0.530 ;
      RECT 0.400 0.595 0.475 1.080 ;
      RECT 0.400 0.175 0.490 0.355 ;
      RECT 0.580 0.345 0.725 0.500 ;
      RECT 0.490 0.175 0.815 0.255 ;
      RECT 0.390 1.145 0.905 1.225 ;
      RECT 0.815 0.175 0.920 0.330 ;
      RECT 0.475 1.010 0.995 1.080 ;
      RECT 0.725 0.420 1.010 0.500 ;
      RECT 0.995 1.010 1.125 1.250 ;
      RECT 1.010 0.295 1.155 0.500 ;
      RECT 1.155 0.295 1.620 0.375 ;
      RECT 1.125 1.035 1.620 1.115 ;
      RECT 1.620 0.295 1.700 1.115 ;
  END
END NCLP3W111OF3X4

MACRO NCLP4W1111OF4X1
  CLASS CORE ;
  FOREIGN NCLP4W1111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.110 0.595 0.665 0.805 ;
        RECT 0.665 0.715 0.960 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.455 0.970 0.530 ;
        RECT 0.970 0.320 1.150 0.530 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.365 0.870 1.145 0.960 ;
        RECT 1.145 0.595 1.235 0.960 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048500 ;
    PORT
      LAYER metal1 ;
        RECT 1.570 0.590 1.890 0.680 ;
        RECT 1.890 0.590 2.100 0.830 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.038500 ;
    PORT
      LAYER metal1 ;
        RECT 2.525 0.245 2.615 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.245 1.485 ;
        RECT 0.245 1.175 0.380 1.485 ;
        RECT 0.380 1.315 0.605 1.485 ;
        RECT 0.605 1.175 0.770 1.485 ;
        RECT 0.770 1.315 2.005 1.485 ;
        RECT 2.005 1.035 2.100 1.485 ;
        RECT 2.100 1.315 2.355 1.485 ;
        RECT 2.355 0.620 2.445 1.485 ;
        RECT 2.445 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.215 0.085 ;
        RECT 0.215 -0.085 0.380 0.255 ;
        RECT 0.380 -0.085 0.605 0.085 ;
        RECT 0.605 -0.085 0.770 0.255 ;
        RECT 0.770 -0.085 1.965 0.085 ;
        RECT 1.965 -0.085 2.060 0.255 ;
        RECT 2.060 -0.085 2.355 0.085 ;
        RECT 2.355 -0.085 2.445 0.450 ;
        RECT 2.445 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.160 0.145 0.390 ;
      RECT 0.045 1.035 0.180 1.240 ;
      RECT 0.145 0.320 0.445 0.390 ;
      RECT 0.445 0.160 0.540 0.390 ;
      RECT 0.540 0.320 0.835 0.390 ;
      RECT 0.835 0.175 0.905 0.390 ;
      RECT 1.300 0.320 1.370 0.970 ;
      RECT 1.435 0.455 1.505 0.815 ;
      RECT 1.370 0.880 1.690 0.970 ;
      RECT 1.505 0.745 1.755 0.815 ;
      RECT 1.755 0.745 1.825 0.970 ;
      RECT 0.905 0.175 1.900 0.255 ;
      RECT 0.180 1.035 1.935 1.110 ;
      RECT 1.370 0.320 2.135 0.390 ;
      RECT 1.825 0.895 2.165 0.970 ;
      RECT 1.505 0.455 2.200 0.525 ;
      RECT 2.200 0.160 2.290 0.525 ;
      RECT 2.165 0.895 2.290 1.195 ;
  END
END NCLP4W1111OF4X1

MACRO NCLP4W1111OF4X2
  CLASS CORE ;
  FOREIGN NCLP4W1111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.090 0.450 0.390 0.670 ;
        RECT 0.390 0.590 0.960 0.670 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.545 0.435 1.170 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.735 0.940 0.805 ;
        RECT 0.940 0.735 1.080 1.085 ;
        RECT 1.080 0.590 1.170 1.085 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050000 ;
    PORT
      LAYER metal1 ;
        RECT 1.370 0.525 1.470 0.825 ;
        RECT 1.470 0.735 1.925 0.825 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079750 ;
    PORT
      LAYER metal1 ;
        RECT 2.165 0.525 2.335 0.645 ;
        RECT 2.335 0.170 2.425 1.210 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.200 1.485 ;
        RECT 0.200 1.005 0.335 1.485 ;
        RECT 0.335 1.315 0.585 1.485 ;
        RECT 0.585 1.005 0.720 1.485 ;
        RECT 0.720 1.315 1.785 1.485 ;
        RECT 1.785 0.945 1.925 1.485 ;
        RECT 1.925 1.315 2.165 1.485 ;
        RECT 2.165 0.710 2.255 1.485 ;
        RECT 2.255 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.200 0.085 ;
        RECT 0.200 -0.085 0.335 0.235 ;
        RECT 0.335 -0.085 0.585 0.085 ;
        RECT 0.585 -0.085 0.720 0.235 ;
        RECT 0.720 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.925 0.245 ;
        RECT 1.925 -0.085 2.165 0.085 ;
        RECT 2.165 -0.085 2.255 0.450 ;
        RECT 2.255 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.170 0.135 0.370 ;
      RECT 0.045 0.870 0.135 1.210 ;
      RECT 0.135 0.300 0.400 0.370 ;
      RECT 0.135 0.870 0.400 0.940 ;
      RECT 0.400 0.170 0.520 0.370 ;
      RECT 0.400 0.870 0.520 1.210 ;
      RECT 0.520 0.300 0.790 0.370 ;
      RECT 0.520 0.870 0.790 0.940 ;
      RECT 0.790 0.870 0.860 1.220 ;
      RECT 0.790 0.175 0.960 0.370 ;
      RECT 1.235 0.310 1.305 0.960 ;
      RECT 1.305 0.890 1.370 0.960 ;
      RECT 1.370 0.890 1.470 1.050 ;
      RECT 0.860 1.150 1.535 1.220 ;
      RECT 1.535 0.450 1.670 0.670 ;
      RECT 0.960 0.175 1.720 0.245 ;
      RECT 1.535 0.945 1.720 1.220 ;
      RECT 1.305 0.310 1.785 0.385 ;
      RECT 1.785 0.310 1.945 0.535 ;
      RECT 1.670 0.600 2.010 0.670 ;
      RECT 2.010 0.170 2.100 1.210 ;
  END
END NCLP4W1111OF4X2

MACRO NCLP4W1111OF4X4
  CLASS CORE ;
  FOREIGN NCLP4W1111OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051500 ;
    PORT
      LAYER metal1 ;
        RECT 0.055 0.455 0.355 0.810 ;
        RECT 0.355 0.730 0.820 0.810 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051500 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.455 1.150 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051500 ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.875 0.915 0.965 ;
        RECT 0.915 0.785 1.195 0.965 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051750 ;
    PORT
      LAYER metal1 ;
        RECT 1.285 0.665 1.540 0.805 ;
        RECT 1.540 0.665 1.840 0.875 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.170500 ;
    PORT
      LAYER metal1 ;
        RECT 2.090 0.515 2.255 1.005 ;
        RECT 2.255 0.515 2.490 0.815 ;
        RECT 2.490 0.515 2.600 1.005 ;
        RECT 2.600 0.350 2.645 1.005 ;
        RECT 2.645 0.350 2.670 0.585 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.220 1.485 ;
        RECT 0.220 1.225 0.355 1.485 ;
        RECT 0.355 1.315 0.610 1.485 ;
        RECT 0.610 1.225 0.780 1.485 ;
        RECT 0.780 1.315 1.820 1.485 ;
        RECT 1.820 1.100 1.910 1.485 ;
        RECT 1.910 1.315 2.310 1.485 ;
        RECT 2.310 1.240 2.485 1.485 ;
        RECT 2.485 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.220 0.085 ;
        RECT 0.220 -0.085 0.355 0.195 ;
        RECT 0.355 -0.085 0.610 0.085 ;
        RECT 0.610 -0.085 0.780 0.195 ;
        RECT 0.780 -0.085 1.900 0.085 ;
        RECT 1.900 -0.085 2.000 0.285 ;
        RECT 2.000 -0.085 2.310 0.085 ;
        RECT 2.310 -0.085 2.400 0.255 ;
        RECT 2.400 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.050 0.180 0.130 0.365 ;
      RECT 0.045 0.990 0.150 1.160 ;
      RECT 0.130 0.285 0.445 0.365 ;
      RECT 0.445 0.180 0.525 0.365 ;
      RECT 1.285 0.430 1.525 0.575 ;
      RECT 0.525 0.285 1.615 0.365 ;
      RECT 1.615 0.285 1.695 0.420 ;
      RECT 0.150 1.080 1.730 1.160 ;
      RECT 1.535 0.150 1.760 0.220 ;
      RECT 1.760 0.150 1.835 0.425 ;
      RECT 1.525 0.505 1.920 0.575 ;
      RECT 1.285 0.940 1.920 1.015 ;
      RECT 1.920 0.505 2.000 1.015 ;
      RECT 1.835 0.350 2.090 0.425 ;
      RECT 2.090 0.180 2.180 0.425 ;
      RECT 2.180 0.345 2.465 0.425 ;
      RECT 2.465 0.180 2.535 0.425 ;
      RECT 2.535 0.180 2.735 0.260 ;
      RECT 2.000 1.095 2.735 1.175 ;
      RECT 2.735 0.180 2.805 1.175 ;
  END
END NCLP4W1111OF4X4

MACRO NCLP4W3111OF4X1
  CLASS CORE ;
  FOREIGN NCLP4W3111OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.550 0.595 0.785 0.945 ;
        RECT 0.785 0.870 2.145 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.850 0.730 1.785 0.805 ;
        RECT 1.785 0.450 1.935 0.805 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.450 1.220 0.665 ;
        RECT 1.220 0.595 1.720 0.665 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047000 ;
    PORT
      LAYER metal1 ;
        RECT 1.285 0.450 1.720 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.080 0.590 2.340 0.665 ;
        RECT 2.340 0.155 2.355 0.665 ;
        RECT 2.355 0.155 2.425 1.155 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.180 1.485 ;
        RECT 0.180 1.010 0.335 1.485 ;
        RECT 0.335 1.315 2.130 1.485 ;
        RECT 2.130 1.145 2.275 1.485 ;
        RECT 2.275 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.180 0.085 ;
        RECT 0.180 -0.085 0.335 0.245 ;
        RECT 0.335 -0.085 1.990 0.085 ;
        RECT 1.990 -0.085 2.275 0.250 ;
        RECT 2.275 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.155 0.115 1.250 ;
      RECT 0.180 0.315 0.270 0.610 ;
      RECT 0.180 0.810 0.400 0.945 ;
      RECT 0.115 0.675 0.445 0.745 ;
      RECT 0.400 0.810 0.470 1.080 ;
      RECT 0.400 0.175 0.900 0.250 ;
      RECT 0.270 0.315 1.005 0.385 ;
      RECT 0.400 1.145 1.275 1.225 ;
      RECT 0.470 1.010 1.340 1.080 ;
      RECT 1.340 1.010 1.465 1.250 ;
      RECT 1.005 0.175 1.475 0.385 ;
      RECT 1.530 1.145 2.065 1.225 ;
      RECT 1.475 0.315 2.080 0.385 ;
      RECT 1.465 1.010 2.210 1.080 ;
      RECT 2.080 0.315 2.275 0.525 ;
      RECT 2.210 0.730 2.290 1.080 ;
  END
END NCLP4W3111OF4X1

MACRO NCLP4W3111OF4X2
  CLASS CORE ;
  FOREIGN NCLP4W3111OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.465 0.540 0.560 0.760 ;
        RECT 0.560 0.540 0.780 0.945 ;
        RECT 0.780 0.875 2.140 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.845 0.735 1.830 0.810 ;
        RECT 1.830 0.585 2.100 0.810 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.595 1.595 0.670 ;
        RECT 1.595 0.450 1.765 0.670 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.450 1.530 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 2.340 0.175 2.425 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.240 1.485 ;
        RECT 0.240 0.975 0.330 1.485 ;
        RECT 0.330 1.315 2.135 1.485 ;
        RECT 2.135 1.145 2.230 1.485 ;
        RECT 2.230 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.330 0.385 ;
        RECT 0.330 -0.085 2.045 0.085 ;
        RECT 2.045 -0.085 2.230 0.385 ;
        RECT 2.230 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.305 0.135 1.250 ;
      RECT 0.205 0.755 0.330 0.910 ;
      RECT 0.135 0.485 0.400 0.690 ;
      RECT 0.330 0.840 0.400 0.910 ;
      RECT 0.400 0.840 0.495 1.080 ;
      RECT 0.400 0.175 0.525 0.420 ;
      RECT 0.590 0.310 0.875 0.475 ;
      RECT 0.525 0.175 0.890 0.245 ;
      RECT 0.875 0.310 1.230 0.385 ;
      RECT 0.395 1.145 1.290 1.225 ;
      RECT 1.230 0.175 1.830 0.385 ;
      RECT 1.830 0.175 1.900 0.520 ;
      RECT 1.525 1.145 2.070 1.225 ;
      RECT 1.900 0.450 2.205 0.520 ;
      RECT 0.495 1.010 2.205 1.080 ;
      RECT 2.205 0.450 2.275 1.080 ;
  END
END NCLP4W3111OF4X2

MACRO NCLPAO22OF4X1
  CLASS CORE ;
  FOREIGN NCLPAO22OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 1.210 0.730 2.080 0.805 ;
        RECT 2.080 0.730 2.320 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.595 1.990 0.665 ;
        RECT 1.990 0.375 2.290 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.720 0.660 1.135 0.945 ;
        RECT 1.135 0.870 1.950 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 1.085 0.445 1.910 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 2.525 0.150 2.615 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.210 1.485 ;
        RECT 0.210 0.660 0.345 1.485 ;
        RECT 0.345 1.315 0.715 1.485 ;
        RECT 0.715 1.145 0.885 1.485 ;
        RECT 0.885 1.315 2.250 1.485 ;
        RECT 2.250 1.225 2.455 1.485 ;
        RECT 2.455 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.210 0.085 ;
        RECT 0.210 -0.085 0.345 0.250 ;
        RECT 0.345 -0.085 2.265 0.085 ;
        RECT 2.265 -0.085 2.455 0.175 ;
        RECT 2.455 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.115 0.910 ;
      RECT 0.115 0.150 0.135 0.460 ;
      RECT 0.135 0.360 0.375 0.460 ;
      RECT 0.440 0.150 0.530 0.460 ;
      RECT 0.440 0.660 0.645 1.080 ;
      RECT 0.595 0.175 0.685 0.325 ;
      RECT 0.530 0.390 0.750 0.460 ;
      RECT 0.750 0.310 0.885 0.460 ;
      RECT 0.180 0.525 0.950 0.595 ;
      RECT 0.645 1.010 0.950 1.080 ;
      RECT 0.950 0.310 1.020 0.595 ;
      RECT 0.950 1.010 1.020 1.225 ;
      RECT 0.685 0.175 1.470 0.245 ;
      RECT 1.020 0.310 1.535 0.380 ;
      RECT 1.535 0.240 1.685 0.380 ;
      RECT 1.020 1.145 1.845 1.225 ;
      RECT 1.685 0.240 2.385 0.310 ;
      RECT 1.100 1.010 2.385 1.080 ;
      RECT 2.385 0.240 2.455 1.080 ;
  END
END NCLPAO22OF4X1

MACRO NCLPAO22OF4X2
  CLASS CORE ;
  FOREIGN NCLPAO22OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 1.260 0.735 2.345 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.595 1.990 0.665 ;
        RECT 1.990 0.420 2.290 0.665 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.810 0.755 1.110 0.945 ;
        RECT 1.110 0.875 2.290 0.945 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.555 0.550 0.720 0.875 ;
        RECT 0.720 0.550 0.850 0.665 ;
        RECT 0.850 0.460 1.150 0.665 ;
        RECT 1.150 0.460 1.730 0.530 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 2.545 0.165 2.615 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 0.975 0.305 1.485 ;
        RECT 0.305 1.315 0.700 1.485 ;
        RECT 0.700 1.290 0.935 1.485 ;
        RECT 0.935 1.315 2.210 1.485 ;
        RECT 2.210 1.170 2.435 1.485 ;
        RECT 2.435 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.225 0.085 ;
        RECT 0.225 -0.085 0.310 0.390 ;
        RECT 0.310 -0.085 2.230 0.085 ;
        RECT 2.230 -0.085 2.450 0.175 ;
        RECT 2.450 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.325 0.115 1.250 ;
      RECT 0.115 0.325 0.135 0.685 ;
      RECT 0.205 0.775 0.395 0.910 ;
      RECT 0.135 0.480 0.435 0.685 ;
      RECT 0.395 0.775 0.465 1.080 ;
      RECT 0.555 0.175 0.690 0.260 ;
      RECT 0.400 0.325 0.750 0.395 ;
      RECT 0.750 0.310 0.885 0.395 ;
      RECT 0.690 0.175 0.950 0.245 ;
      RECT 0.950 0.175 1.450 0.260 ;
      RECT 1.095 0.325 1.540 0.395 ;
      RECT 1.540 0.260 1.650 0.395 ;
      RECT 0.395 1.145 1.835 1.215 ;
      RECT 1.650 0.260 2.410 0.330 ;
      RECT 0.465 1.010 2.410 1.080 ;
      RECT 2.410 0.260 2.480 1.080 ;
  END
END NCLPAO22OF4X2

MACRO NCLPOA22OF4X1
  CLASS CORE ;
  FOREIGN NCLPOA22OF4X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.870 1.890 0.945 ;
        RECT 1.890 0.590 2.100 0.945 ;
        RECT 2.100 0.590 2.320 0.805 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 0.710 0.455 0.975 0.805 ;
        RECT 0.975 0.455 2.160 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.590 1.805 0.670 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 1.040 0.735 1.720 0.805 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 2.525 0.155 2.615 1.245 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.200 1.485 ;
        RECT 0.200 0.730 0.335 1.485 ;
        RECT 0.335 1.315 1.830 1.485 ;
        RECT 1.830 1.280 2.040 1.485 ;
        RECT 2.040 1.315 2.325 1.485 ;
        RECT 2.325 1.145 2.460 1.485 ;
        RECT 2.460 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.335 0.255 ;
        RECT 0.335 -0.085 2.190 0.085 ;
        RECT 2.190 -0.085 2.405 0.220 ;
        RECT 2.405 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.155 0.120 0.975 ;
      RECT 0.120 0.455 0.135 0.975 ;
      RECT 0.135 0.455 0.445 0.665 ;
      RECT 0.425 0.730 0.495 1.225 ;
      RECT 0.415 0.175 1.110 0.255 ;
      RECT 0.185 0.320 1.275 0.390 ;
      RECT 0.495 1.145 1.290 1.225 ;
      RECT 1.485 1.145 2.260 1.215 ;
      RECT 1.275 0.300 2.385 0.390 ;
      RECT 0.560 1.010 2.385 1.080 ;
      RECT 2.385 0.300 2.460 1.080 ;
  END
END NCLPOA22OF4X1

MACRO NCLPOA22OF4X2
  CLASS CORE ;
  FOREIGN NCLPOA22OF4X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.635 0.730 0.945 ;
        RECT 0.730 0.875 2.150 0.945 ;
        RECT 2.150 0.635 2.290 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.820 0.455 1.035 0.735 ;
        RECT 1.035 0.455 2.290 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.595 1.945 0.670 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 1.125 0.735 1.910 0.805 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078650 ;
    PORT
      LAYER metal1 ;
        RECT 2.545 0.160 2.615 1.225 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.225 1.485 ;
        RECT 0.225 0.865 0.320 1.485 ;
        RECT 0.320 1.315 1.910 1.485 ;
        RECT 1.910 1.290 2.045 1.485 ;
        RECT 2.045 1.315 2.355 1.485 ;
        RECT 2.355 1.150 2.445 1.485 ;
        RECT 2.445 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.205 0.085 ;
        RECT 0.205 -0.085 0.320 0.240 ;
        RECT 0.320 -0.085 2.290 0.085 ;
        RECT 2.290 -0.085 2.395 0.230 ;
        RECT 2.395 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.115 1.140 ;
      RECT 0.115 0.570 0.135 1.140 ;
      RECT 0.135 0.570 0.475 0.775 ;
      RECT 0.410 0.865 0.500 1.225 ;
      RECT 0.205 0.320 0.710 0.480 ;
      RECT 0.410 0.175 1.155 0.250 ;
      RECT 0.500 1.155 1.330 1.225 ;
      RECT 0.710 0.320 1.365 0.390 ;
      RECT 1.365 0.230 1.515 0.390 ;
      RECT 1.555 1.145 2.265 1.215 ;
      RECT 1.515 0.320 2.385 0.390 ;
      RECT 0.565 1.010 2.385 1.080 ;
      RECT 2.385 0.320 2.460 1.080 ;
  END
END NCLPOA22OF4X2

MACRO NCLPOA22OF4X4
  CLASS CORE ;
  FOREIGN NCLPOA22OF4X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.850 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.665 0.715 0.800 0.945 ;
        RECT 0.800 0.875 2.130 0.945 ;
        RECT 2.130 0.650 2.265 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.890 0.455 1.025 0.715 ;
        RECT 1.025 0.455 2.170 0.525 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.590 1.940 0.665 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 1.115 0.730 1.720 0.810 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105850 ;
    PORT
      LAYER metal1 ;
        RECT 2.530 0.175 2.620 1.235 ;
        RECT 2.620 0.500 2.790 0.760 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.205 1.485 ;
        RECT 0.205 0.740 0.340 1.485 ;
        RECT 0.340 1.315 1.855 1.485 ;
        RECT 1.855 1.290 2.035 1.485 ;
        RECT 2.035 1.315 2.345 1.485 ;
        RECT 2.345 1.170 2.435 1.485 ;
        RECT 2.435 1.315 2.715 1.485 ;
        RECT 2.715 0.890 2.805 1.485 ;
        RECT 2.805 1.315 2.850 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.240 0.085 ;
        RECT 0.240 -0.085 0.330 0.255 ;
        RECT 0.330 -0.085 2.270 0.085 ;
        RECT 2.270 -0.085 2.450 0.210 ;
        RECT 2.450 -0.085 2.715 0.085 ;
        RECT 2.715 -0.085 2.805 0.390 ;
        RECT 2.805 -0.085 2.850 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.210 0.125 0.980 ;
      RECT 0.430 0.740 0.500 1.225 ;
      RECT 0.125 0.570 0.585 0.650 ;
      RECT 0.205 0.345 0.610 0.480 ;
      RECT 0.610 0.320 0.750 0.480 ;
      RECT 0.420 0.175 1.110 0.255 ;
      RECT 0.750 0.320 1.300 0.390 ;
      RECT 0.500 1.145 1.300 1.225 ;
      RECT 1.510 1.145 2.255 1.225 ;
      RECT 1.300 0.300 2.360 0.390 ;
      RECT 0.565 1.010 2.360 1.080 ;
      RECT 2.360 0.300 2.450 1.080 ;
  END
END NCLPOA22OF4X4

MACRO PULLDOWN
  CLASS CORE TIELOW ;
  FOREIGN PULLDOWN 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.380 BY 1.400 ;
  PIN Q
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.032450 ;
    ANTENNAGATEAREA 0.014750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.435 0.245 0.735 ;
        RECT 0.245 0.150 0.335 0.735 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.380 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.075 0.085 ;
        RECT 0.075 -0.085 0.175 0.355 ;
        RECT 0.175 -0.085 0.380 0.085 ;
    END
  END VSS
END PULLDOWN

MACRO PULLUP
  CLASS CORE TIEHIGH ;
  FOREIGN PULLUP 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 0.380 BY 1.400 ;
  PIN Q
    DIRECTION INOUT ;
    ANTENNADIFFAREA 0.044550 ;
    ANTENNAGATEAREA 0.020250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.525 0.245 0.810 ;
        RECT 0.245 0.525 0.335 1.250 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.075 1.485 ;
        RECT 0.075 0.875 0.165 1.485 ;
        RECT 0.165 1.315 0.380 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.380 0.085 ;
    END
  END VSS
END PULLUP

MACRO RACELEM1X1
  CLASS CORE ;
  FOREIGN RACELEM1X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.340 0.810 0.420 0.945 ;
        RECT 0.420 0.870 0.960 0.945 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022750 ;
    PORT
      LAYER metal1 ;
        RECT 0.630 0.355 1.080 0.595 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.024750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.525 0.130 0.940 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.034100 ;
    PORT
      LAYER metal1 ;
        RECT 1.955 0.245 2.045 1.015 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.505 0.685 0.750 0.765 ;
        RECT 0.750 0.685 1.080 0.805 ;
        RECT 1.080 0.685 1.380 0.945 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.030 0.125 1.485 ;
        RECT 0.125 1.315 1.235 1.485 ;
        RECT 1.235 1.170 1.345 1.485 ;
        RECT 1.345 1.315 1.785 1.485 ;
        RECT 1.785 0.675 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.890 0.085 ;
        RECT 0.890 -0.085 1.145 0.110 ;
        RECT 1.145 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.865 0.545 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.450 ;
      RECT 0.125 0.350 0.205 0.450 ;
      RECT 0.205 0.350 0.275 1.080 ;
      RECT 0.275 0.350 0.540 0.440 ;
      RECT 0.505 1.145 1.145 1.225 ;
      RECT 0.275 1.010 1.435 1.080 ;
      RECT 1.435 1.010 1.445 1.250 ;
      RECT 1.445 0.575 1.525 1.250 ;
      RECT 1.525 0.575 1.560 0.710 ;
      RECT 1.160 0.355 1.625 0.490 ;
      RECT 1.590 0.800 1.625 0.945 ;
      RECT 1.625 0.355 1.695 0.945 ;
      RECT 0.215 0.185 1.700 0.265 ;
  END
END RACELEM1X1

MACRO RACELEM1X2
  CLASS CORE ;
  FOREIGN RACELEM1X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.735 0.960 0.825 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.021750 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.435 1.025 0.525 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.525 0.130 0.875 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.075600 ;
    PORT
      LAYER metal1 ;
        RECT 1.955 0.240 2.045 1.165 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.490 0.590 1.145 0.670 ;
        RECT 1.145 0.590 1.400 0.875 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.965 0.125 1.485 ;
        RECT 0.125 1.315 1.210 1.485 ;
        RECT 1.210 1.135 1.345 1.485 ;
        RECT 1.345 1.315 1.775 1.485 ;
        RECT 1.775 0.950 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.950 0.085 ;
        RECT 0.950 -0.085 1.130 0.165 ;
        RECT 1.130 -0.085 1.775 0.085 ;
        RECT 1.775 -0.085 1.865 0.475 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 0.460 ;
      RECT 0.125 0.380 0.215 0.460 ;
      RECT 0.215 0.380 0.290 1.045 ;
      RECT 0.205 0.175 0.340 0.285 ;
      RECT 0.290 0.965 0.400 1.045 ;
      RECT 0.290 0.380 0.410 0.475 ;
      RECT 0.410 0.335 0.490 0.475 ;
      RECT 0.400 0.965 0.490 1.225 ;
      RECT 0.340 0.175 0.610 0.245 ;
      RECT 0.610 0.175 0.690 0.330 ;
      RECT 0.580 1.135 1.125 1.225 ;
      RECT 0.490 0.965 1.435 1.045 ;
      RECT 1.435 0.965 1.465 1.225 ;
      RECT 1.465 0.590 1.540 1.225 ;
      RECT 1.095 0.420 1.605 0.500 ;
      RECT 0.690 0.250 1.665 0.330 ;
      RECT 1.605 0.420 1.685 1.225 ;
  END
END RACELEM1X2

MACRO RACELEM1X4
  CLASS CORE ;
  FOREIGN RACELEM1X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.355 0.735 0.605 0.945 ;
        RECT 0.605 0.855 0.770 0.945 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.315 1.015 0.525 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.510 0.130 0.785 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.103675 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.235 2.050 1.240 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.435 0.590 0.860 0.670 ;
        RECT 0.860 0.590 0.945 0.920 ;
        RECT 0.945 0.645 1.330 0.920 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.995 0.125 1.485 ;
        RECT 0.125 1.315 1.195 1.485 ;
        RECT 1.195 1.170 1.330 1.485 ;
        RECT 1.330 1.315 1.770 1.485 ;
        RECT 1.770 0.965 1.870 1.485 ;
        RECT 1.870 1.315 2.145 1.485 ;
        RECT 2.145 0.885 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.915 0.085 ;
        RECT 0.915 -0.085 1.120 0.110 ;
        RECT 1.120 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.870 0.420 ;
        RECT 1.870 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.445 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.150 0.125 0.425 ;
      RECT 0.125 0.345 0.215 0.425 ;
      RECT 0.215 0.345 0.290 1.080 ;
      RECT 0.290 0.345 0.390 0.425 ;
      RECT 0.390 0.325 0.530 0.425 ;
      RECT 0.540 1.145 1.120 1.225 ;
      RECT 0.290 1.010 1.420 1.080 ;
      RECT 1.420 0.645 1.500 1.235 ;
      RECT 0.205 0.175 1.535 0.250 ;
      RECT 1.590 0.815 1.680 1.100 ;
      RECT 1.105 0.395 1.705 0.555 ;
      RECT 1.500 0.645 1.710 0.725 ;
      RECT 1.705 0.485 1.790 0.555 ;
      RECT 1.680 0.815 1.790 0.895 ;
      RECT 1.790 0.485 1.870 0.895 ;
  END
END RACELEM1X4

MACRO RACELEM2X1
  CLASS CORE ;
  FOREIGN RACELEM2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.053000 ;
    PORT
      LAYER metal1 ;
        RECT 0.525 0.595 0.660 0.825 ;
        RECT 0.660 0.595 1.530 0.670 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022750 ;
    PORT
      LAYER metal1 ;
        RECT 0.130 0.595 0.390 0.825 ;
    END
  END M1
  PIN M2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.022750 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.310 0.370 0.530 ;
        RECT 0.370 0.220 0.460 0.530 ;
    END
  END M2
  PIN P1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.030250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.450 1.035 0.530 ;
    END
  END P1
  PIN P2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.030250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.450 1.530 0.530 ;
    END
  END P2
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.035700 ;
    PORT
      LAYER metal1 ;
        RECT 2.340 0.220 2.425 1.155 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.056000 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.735 1.565 0.825 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.820 1.485 ;
        RECT 0.820 1.240 1.035 1.485 ;
        RECT 1.035 1.315 1.820 1.485 ;
        RECT 1.820 0.975 1.920 1.485 ;
        RECT 1.920 1.315 2.170 1.485 ;
        RECT 2.170 0.645 2.250 1.485 ;
        RECT 2.250 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.115 0.405 ;
        RECT 0.115 -0.085 1.805 0.085 ;
        RECT 1.805 -0.085 1.895 0.390 ;
        RECT 1.895 -0.085 2.170 0.085 ;
        RECT 2.170 -0.085 2.250 0.440 ;
        RECT 2.250 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.915 0.145 1.170 ;
      RECT 0.820 0.220 0.920 0.380 ;
      RECT 1.010 0.175 1.565 0.245 ;
      RECT 0.920 0.310 1.635 0.380 ;
      RECT 0.235 0.920 1.635 1.010 ;
      RECT 1.635 0.310 1.715 1.010 ;
      RECT 0.145 1.090 1.725 1.170 ;
      RECT 1.715 0.480 1.920 0.615 ;
      RECT 1.805 0.680 1.985 0.885 ;
      RECT 1.985 0.310 2.080 0.885 ;
  END
END RACELEM2X1

MACRO RACELEM2X2
  CLASS CORE ;
  FOREIGN RACELEM2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.053750 ;
    PORT
      LAYER metal1 ;
        RECT 0.505 0.595 1.530 0.670 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025000 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.595 0.390 0.875 ;
    END
  END M1
  PIN M2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.175 0.460 0.525 ;
    END
  END M2
  PIN P1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.028750 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.450 1.020 0.530 ;
    END
  END P1
  PIN P2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.028750 ;
    PORT
      LAYER metal1 ;
        RECT 1.110 0.450 1.720 0.530 ;
    END
  END P2
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.078650 ;
    PORT
      LAYER metal1 ;
        RECT 2.335 0.150 2.425 1.160 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.055000 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.735 1.620 0.825 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.795 1.485 ;
        RECT 0.795 1.240 0.960 1.485 ;
        RECT 0.960 1.315 1.800 1.485 ;
        RECT 1.800 1.105 1.885 1.485 ;
        RECT 1.885 1.315 2.155 1.485 ;
        RECT 2.155 0.760 2.245 1.485 ;
        RECT 2.245 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.115 0.415 ;
        RECT 0.115 -0.085 1.695 0.085 ;
        RECT 1.695 -0.085 1.915 0.220 ;
        RECT 1.915 -0.085 2.155 0.085 ;
        RECT 2.155 -0.085 2.245 0.220 ;
        RECT 2.245 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.965 0.125 1.240 ;
      RECT 0.125 1.080 0.185 1.240 ;
      RECT 0.795 0.175 0.935 0.380 ;
      RECT 1.005 0.175 1.530 0.245 ;
      RECT 0.185 1.080 1.710 1.160 ;
      RECT 0.935 0.310 1.785 0.380 ;
      RECT 0.210 0.940 1.785 1.015 ;
      RECT 1.785 0.310 1.865 1.015 ;
      RECT 1.865 0.310 1.915 0.555 ;
      RECT 1.935 0.645 1.975 0.940 ;
      RECT 1.975 0.645 1.980 1.200 ;
      RECT 1.980 0.175 2.065 1.200 ;
  END
END RACELEM2X2

MACRO RACELEM2X4
  CLASS CORE ;
  FOREIGN RACELEM2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.051500 ;
    PORT
      LAYER metal1 ;
        RECT 0.510 0.595 0.660 0.860 ;
        RECT 0.660 0.595 1.530 0.670 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.595 0.390 0.875 ;
    END
  END M1
  PIN M2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.250 0.175 0.580 0.505 ;
    END
  END M2
  PIN P1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.027750 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.450 1.040 0.530 ;
    END
  END P1
  PIN P2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.027750 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.450 1.340 0.530 ;
    END
  END P2
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 2.175 0.625 2.335 0.715 ;
        RECT 2.335 0.150 2.425 1.030 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER metal1 ;
        RECT 0.750 0.735 1.560 0.825 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.800 1.485 ;
        RECT 0.800 1.240 0.990 1.485 ;
        RECT 0.990 1.315 1.795 1.485 ;
        RECT 1.795 0.975 1.875 1.485 ;
        RECT 1.875 1.315 2.155 1.485 ;
        RECT 2.155 0.805 2.245 1.485 ;
        RECT 2.245 1.315 2.525 1.485 ;
        RECT 2.525 0.805 2.615 1.485 ;
        RECT 2.615 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.060 0.085 ;
        RECT 0.060 -0.085 0.160 0.410 ;
        RECT 0.160 -0.085 1.775 0.085 ;
        RECT 1.775 -0.085 1.910 0.380 ;
        RECT 1.910 -0.085 2.155 0.085 ;
        RECT 2.155 -0.085 2.245 0.505 ;
        RECT 2.245 -0.085 2.525 0.085 ;
        RECT 2.525 -0.085 2.615 0.505 ;
        RECT 2.615 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.965 0.125 1.240 ;
      RECT 0.125 1.095 0.215 1.240 ;
      RECT 0.800 0.175 0.935 0.385 ;
      RECT 0.935 0.315 1.430 0.385 ;
      RECT 1.430 0.315 1.510 0.505 ;
      RECT 1.005 0.175 1.555 0.250 ;
      RECT 1.510 0.425 1.625 0.505 ;
      RECT 0.215 0.950 1.625 1.030 ;
      RECT 1.625 0.425 1.700 1.030 ;
      RECT 1.700 0.635 1.705 1.030 ;
      RECT 0.215 1.095 1.715 1.175 ;
      RECT 1.790 0.805 1.965 0.885 ;
      RECT 1.790 0.465 2.065 0.545 ;
      RECT 1.965 0.805 2.065 1.080 ;
      RECT 1.705 0.635 2.085 0.715 ;
  END
END RACELEM2X4

MACRO RNCL2W11OF2X1
  CLASS CORE ;
  FOREIGN RNCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.845 0.870 1.575 0.950 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.455 1.175 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.225 2.045 1.230 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.045500 ;
    PORT
      LAYER metal1 ;
        RECT 0.550 0.730 0.755 0.900 ;
        RECT 0.755 0.730 1.760 0.805 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.215 1.485 ;
        RECT 0.215 0.945 0.295 1.485 ;
        RECT 0.295 1.315 0.735 1.485 ;
        RECT 0.735 1.290 0.920 1.485 ;
        RECT 0.920 1.315 1.785 1.485 ;
        RECT 1.785 1.085 1.870 1.485 ;
        RECT 1.870 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.235 0.085 ;
        RECT 0.235 -0.085 0.390 0.310 ;
        RECT 0.390 -0.085 1.630 0.085 ;
        RECT 1.630 -0.085 1.850 0.245 ;
        RECT 1.850 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.225 0.125 1.220 ;
      RECT 0.125 0.650 0.460 0.855 ;
      RECT 0.385 0.970 0.485 1.225 ;
      RECT 0.195 0.410 0.735 0.560 ;
      RECT 0.735 0.320 0.845 0.560 ;
      RECT 0.575 0.175 1.065 0.255 ;
      RECT 0.845 0.320 1.145 0.390 ;
      RECT 1.145 0.180 1.280 0.390 ;
      RECT 0.485 1.150 1.470 1.225 ;
      RECT 0.575 1.015 1.555 1.085 ;
      RECT 1.555 1.015 1.640 1.225 ;
      RECT 1.640 0.915 1.720 1.225 ;
      RECT 1.280 0.310 1.825 0.390 ;
      RECT 1.720 0.915 1.825 0.995 ;
      RECT 1.825 0.310 1.895 0.995 ;
  END
END RNCL2W11OF2X1

MACRO RNCL2W11OF2X2
  CLASS CORE ;
  FOREIGN RNCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.835 0.735 1.545 0.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.047500 ;
    PORT
      LAYER metal1 ;
        RECT 0.940 0.455 1.200 0.530 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.230 2.045 1.220 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.046500 ;
    PORT
      LAYER metal1 ;
        RECT 0.540 0.595 0.745 0.815 ;
        RECT 0.745 0.595 1.760 0.670 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.230 1.485 ;
        RECT 0.230 0.880 0.320 1.485 ;
        RECT 0.320 1.315 0.745 1.485 ;
        RECT 0.745 1.180 0.880 1.485 ;
        RECT 0.880 1.315 1.715 1.485 ;
        RECT 1.715 1.150 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.230 0.085 ;
        RECT 0.230 -0.085 0.450 0.220 ;
        RECT 0.450 -0.085 1.665 0.085 ;
        RECT 1.665 -0.085 1.850 0.380 ;
        RECT 1.850 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.175 0.125 1.155 ;
      RECT 0.125 0.585 0.135 1.155 ;
      RECT 0.205 0.310 0.405 0.495 ;
      RECT 0.135 0.585 0.450 0.790 ;
      RECT 0.410 0.905 0.500 1.225 ;
      RECT 0.500 1.045 0.560 1.225 ;
      RECT 0.560 1.045 0.970 1.115 ;
      RECT 0.970 1.045 1.050 1.225 ;
      RECT 0.590 0.175 1.075 0.245 ;
      RECT 0.590 0.905 1.140 0.980 ;
      RECT 0.405 0.310 1.145 0.390 ;
      RECT 1.145 0.175 1.350 0.390 ;
      RECT 1.350 0.175 1.430 0.525 ;
      RECT 1.050 1.150 1.465 1.225 ;
      RECT 1.430 0.445 1.825 0.525 ;
      RECT 1.140 0.905 1.825 1.060 ;
      RECT 1.825 0.445 1.895 1.060 ;
  END
END RNCL2W11OF2X2

MACRO RNCL2W11OF2X4
  CLASS CORE ;
  FOREIGN RNCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.058500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.640 0.510 0.875 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.058500 ;
    PORT
      LAYER metal1 ;
        RECT 0.090 0.455 0.660 0.545 ;
        RECT 0.660 0.455 0.960 0.705 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.103675 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.175 2.050 1.170 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.028250 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.455 1.650 0.735 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 0.970 0.125 1.485 ;
        RECT 0.125 1.315 0.385 1.485 ;
        RECT 0.385 1.100 0.535 1.485 ;
        RECT 0.535 1.315 1.390 1.485 ;
        RECT 1.390 0.990 1.495 1.485 ;
        RECT 1.495 1.315 1.745 1.485 ;
        RECT 1.745 0.985 1.880 1.485 ;
        RECT 1.880 1.315 2.145 1.485 ;
        RECT 2.145 0.810 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.380 ;
        RECT 0.125 -0.085 0.385 0.085 ;
        RECT 0.385 -0.085 0.535 0.220 ;
        RECT 0.535 -0.085 1.715 0.085 ;
        RECT 1.715 -0.085 1.880 0.110 ;
        RECT 1.880 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.375 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 0.950 0.295 1.225 ;
      RECT 0.295 0.950 0.875 1.030 ;
      RECT 0.875 0.950 1.000 1.225 ;
      RECT 0.720 0.795 1.050 0.875 ;
      RECT 1.050 0.460 1.065 0.875 ;
      RECT 0.200 0.310 1.075 0.380 ;
      RECT 1.065 0.460 1.135 1.095 ;
      RECT 1.135 0.460 1.165 0.545 ;
      RECT 1.135 1.015 1.165 1.095 ;
      RECT 1.165 0.320 1.245 0.545 ;
      RECT 1.200 0.790 1.280 0.925 ;
      RECT 0.720 0.175 1.300 0.245 ;
      RECT 1.165 1.015 1.300 1.225 ;
      RECT 1.280 0.845 1.585 0.925 ;
      RECT 1.585 0.845 1.600 1.225 ;
      RECT 1.245 0.320 1.620 0.390 ;
      RECT 1.600 0.800 1.665 1.225 ;
      RECT 1.505 0.175 1.745 0.255 ;
      RECT 1.665 0.800 1.745 0.895 ;
      RECT 1.745 0.175 1.825 0.895 ;
  END
END RNCL2W11OF2X4

MACRO RSNCL2W11OF2X1
  CLASS CORE ;
  FOREIGN RSNCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.550 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.855 0.640 0.945 ;
        RECT 0.640 0.600 0.795 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040700 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.765 2.145 0.855 ;
        RECT 2.145 0.245 2.235 1.220 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.315 1.570 0.450 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 1.110 0.525 1.315 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.125 1.485 ;
        RECT 0.125 1.315 0.430 1.485 ;
        RECT 0.430 1.180 0.550 1.485 ;
        RECT 0.550 1.315 1.530 1.485 ;
        RECT 1.530 1.290 1.715 1.485 ;
        RECT 1.715 1.315 1.960 1.485 ;
        RECT 1.960 0.945 2.050 1.485 ;
        RECT 2.050 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.435 ;
        RECT 0.130 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.550 0.265 ;
        RECT 0.550 -0.085 1.110 0.085 ;
        RECT 1.110 -0.085 1.265 0.110 ;
        RECT 1.265 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.050 0.455 ;
        RECT 2.050 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.160 0.310 0.435 ;
      RECT 0.205 1.010 0.340 1.225 ;
      RECT 0.340 1.010 0.900 1.090 ;
      RECT 0.715 0.175 0.915 0.265 ;
      RECT 0.310 0.355 0.975 0.435 ;
      RECT 0.900 0.955 1.070 1.090 ;
      RECT 0.975 0.335 1.110 0.435 ;
      RECT 0.700 1.155 1.135 1.225 ;
      RECT 1.135 1.065 1.205 1.225 ;
      RECT 0.885 0.800 1.270 0.880 ;
      RECT 1.270 0.800 1.340 1.220 ;
      RECT 0.915 0.175 1.495 0.250 ;
      RECT 1.405 0.690 1.495 1.010 ;
      RECT 1.340 1.100 1.585 1.220 ;
      RECT 1.495 0.690 1.635 0.795 ;
      RECT 1.635 0.175 1.715 0.795 ;
      RECT 1.585 0.980 1.780 1.220 ;
      RECT 1.780 0.400 1.870 1.220 ;
  END
END RSNCL2W11OF2X1

MACRO RSNCL2W11OF2X2
  CLASS CORE ;
  FOREIGN RSNCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.053000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.550 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.053000 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.855 0.640 0.945 ;
        RECT 0.640 0.600 0.795 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.080300 ;
    PORT
      LAYER metal1 ;
        RECT 2.095 0.715 2.145 1.015 ;
        RECT 2.145 0.245 2.235 1.015 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.315 1.570 0.450 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 1.110 0.525 1.315 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.125 1.485 ;
        RECT 0.125 1.315 0.430 1.485 ;
        RECT 0.430 1.180 0.520 1.485 ;
        RECT 0.520 1.315 1.530 1.485 ;
        RECT 1.530 1.275 1.715 1.485 ;
        RECT 1.715 1.315 1.950 1.485 ;
        RECT 1.950 1.090 2.040 1.485 ;
        RECT 2.040 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.415 ;
        RECT 0.125 -0.085 0.430 0.085 ;
        RECT 0.430 -0.085 0.520 0.275 ;
        RECT 0.520 -0.085 1.105 0.085 ;
        RECT 1.105 -0.085 1.265 0.110 ;
        RECT 1.265 -0.085 1.950 0.085 ;
        RECT 1.950 -0.085 2.040 0.495 ;
        RECT 2.040 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.205 0.175 0.340 0.435 ;
      RECT 0.205 1.010 0.340 1.225 ;
      RECT 0.715 0.175 0.880 0.275 ;
      RECT 0.340 1.010 0.900 1.090 ;
      RECT 0.340 0.365 0.970 0.435 ;
      RECT 0.900 0.955 1.070 1.090 ;
      RECT 0.970 0.315 1.110 0.435 ;
      RECT 0.700 1.155 1.135 1.225 ;
      RECT 1.135 1.065 1.205 1.225 ;
      RECT 0.885 0.800 1.270 0.880 ;
      RECT 1.270 0.800 1.340 1.185 ;
      RECT 0.880 0.175 1.495 0.245 ;
      RECT 1.405 0.715 1.495 0.995 ;
      RECT 1.495 0.715 1.635 0.825 ;
      RECT 1.635 0.190 1.715 0.825 ;
      RECT 1.340 1.085 1.780 1.185 ;
      RECT 1.780 0.400 1.860 1.185 ;
  END
END RSNCL2W11OF2X2

MACRO RSNCL2W11OF2X4
  CLASS CORE ;
  FOREIGN RSNCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.585 0.580 0.665 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.735 0.815 0.825 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.104400 ;
    PORT
      LAYER metal1 ;
        RECT 2.145 0.225 2.235 1.155 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 1.390 0.385 1.520 0.660 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 1.200 0.385 1.300 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.000 0.135 1.485 ;
        RECT 0.135 1.315 0.405 1.485 ;
        RECT 0.405 1.160 0.525 1.485 ;
        RECT 0.525 1.315 1.580 1.485 ;
        RECT 1.580 1.260 1.715 1.485 ;
        RECT 1.715 1.315 1.960 1.485 ;
        RECT 1.960 0.895 2.055 1.485 ;
        RECT 2.055 1.315 2.335 1.485 ;
        RECT 2.335 0.755 2.425 1.485 ;
        RECT 2.425 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.495 ;
        RECT 0.130 -0.085 0.390 0.085 ;
        RECT 0.390 -0.085 0.525 0.325 ;
        RECT 0.525 -0.085 1.175 0.085 ;
        RECT 1.175 -0.085 1.310 0.160 ;
        RECT 1.310 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.055 0.455 ;
        RECT 2.055 -0.085 2.335 0.085 ;
        RECT 2.335 -0.085 2.425 0.455 ;
        RECT 2.425 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.220 0.300 0.495 ;
      RECT 0.225 0.935 0.315 1.225 ;
      RECT 0.735 0.225 0.900 0.325 ;
      RECT 0.300 0.415 0.960 0.495 ;
      RECT 0.315 0.935 1.055 1.070 ;
      RECT 0.960 0.395 1.095 0.495 ;
      RECT 0.905 0.710 1.110 0.870 ;
      RECT 0.755 1.145 1.130 1.225 ;
      RECT 1.130 0.950 1.210 1.225 ;
      RECT 1.110 0.800 1.275 0.870 ;
      RECT 1.275 0.800 1.345 1.170 ;
      RECT 0.900 0.225 1.505 0.305 ;
      RECT 1.410 0.865 1.610 1.000 ;
      RECT 1.610 0.190 1.700 1.000 ;
      RECT 1.345 1.090 1.780 1.170 ;
      RECT 1.780 0.395 1.870 1.170 ;
  END
END RSNCL2W11OF2X4

MACRO SACELEM1X1
  CLASS CORE ;
  FOREIGN SACELEM1X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.595 0.580 0.945 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023250 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.130 0.695 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 0.675 0.525 1.080 0.805 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.036300 ;
    PORT
      LAYER metal1 ;
        RECT 1.770 0.495 1.955 0.575 ;
        RECT 1.955 0.310 2.045 0.940 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.048750 ;
    PORT
      LAYER metal1 ;
        RECT 0.815 0.870 1.535 0.955 ;
        RECT 1.535 0.870 1.625 0.995 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.880 1.485 ;
        RECT 0.880 1.215 1.100 1.485 ;
        RECT 1.100 1.315 1.770 1.485 ;
        RECT 1.770 0.665 1.860 1.485 ;
        RECT 1.860 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.295 ;
        RECT 0.125 -0.085 1.195 0.085 ;
        RECT 1.195 -0.085 1.330 0.270 ;
        RECT 1.330 -0.085 1.770 0.085 ;
        RECT 1.770 -0.085 1.860 0.405 ;
        RECT 1.860 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.960 0.125 1.235 ;
      RECT 0.125 0.960 0.210 1.080 ;
      RECT 0.210 0.160 0.280 1.080 ;
      RECT 0.280 0.160 0.490 0.435 ;
      RECT 0.280 1.010 0.545 1.080 ;
      RECT 0.205 1.145 0.710 1.225 ;
      RECT 0.710 1.045 0.790 1.225 ;
      RECT 0.490 0.345 0.910 0.435 ;
      RECT 0.580 0.180 1.110 0.270 ;
      RECT 0.790 1.045 1.190 1.125 ;
      RECT 0.910 0.360 1.315 0.435 ;
      RECT 1.315 0.360 1.420 0.600 ;
      RECT 1.190 1.045 1.455 1.215 ;
      RECT 1.420 0.170 1.525 0.600 ;
      RECT 1.160 0.690 1.590 0.780 ;
      RECT 1.590 0.340 1.680 0.780 ;
  END
END SACELEM1X1

MACRO SACELEM1X2
  CLASS CORE ;
  FOREIGN SACELEM1X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.050250 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.455 0.580 0.805 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.130 0.695 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026500 ;
    PORT
      LAYER metal1 ;
        RECT 0.720 0.665 1.080 0.955 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.785 0.320 1.955 0.620 ;
        RECT 1.955 0.175 2.045 1.060 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.870 0.455 1.180 0.545 ;
        RECT 1.180 0.455 1.375 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.975 1.485 ;
        RECT 0.975 1.215 1.115 1.485 ;
        RECT 1.115 1.315 1.785 1.485 ;
        RECT 1.785 0.845 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.295 ;
        RECT 0.125 -0.085 1.180 0.085 ;
        RECT 1.180 -0.085 1.315 0.240 ;
        RECT 1.315 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.865 0.245 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.820 0.125 1.225 ;
      RECT 0.125 0.820 0.210 0.955 ;
      RECT 0.210 0.310 0.280 0.955 ;
      RECT 0.205 1.020 0.345 1.225 ;
      RECT 0.280 0.310 0.395 0.390 ;
      RECT 0.280 0.875 0.435 0.955 ;
      RECT 0.395 0.175 0.530 0.390 ;
      RECT 0.435 0.875 0.555 1.075 ;
      RECT 0.345 1.145 0.805 1.225 ;
      RECT 0.805 1.045 0.885 1.225 ;
      RECT 0.595 0.175 1.115 0.250 ;
      RECT 0.530 0.315 1.390 0.390 ;
      RECT 1.390 0.175 1.445 0.390 ;
      RECT 0.885 1.045 1.500 1.125 ;
      RECT 1.445 0.175 1.525 0.695 ;
      RECT 1.170 0.820 1.590 0.955 ;
      RECT 1.590 0.175 1.615 0.310 ;
      RECT 1.590 0.820 1.615 1.120 ;
      RECT 1.615 0.175 1.695 1.120 ;
  END
END SACELEM1X2

MACRO SACELEM1X4
  CLASS CORE ;
  FOREIGN SACELEM1X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049750 ;
    PORT
      LAYER metal1 ;
        RECT 0.370 0.455 0.580 0.805 ;
    END
  END A
  PIN M
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.023750 ;
    PORT
      LAYER metal1 ;
        RECT 0.045 0.385 0.130 0.735 ;
    END
  END M
  PIN P
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.720 0.595 0.960 0.945 ;
    END
  END P
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105850 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.245 2.050 1.170 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049250 ;
    PORT
      LAYER metal1 ;
        RECT 0.860 0.455 1.145 0.530 ;
        RECT 1.145 0.455 1.375 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.950 1.485 ;
        RECT 0.950 1.205 1.125 1.485 ;
        RECT 1.125 1.315 1.780 1.485 ;
        RECT 1.780 0.700 1.870 1.485 ;
        RECT 1.870 1.315 2.145 1.485 ;
        RECT 2.145 0.770 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.280 ;
        RECT 0.125 -0.085 1.215 0.085 ;
        RECT 1.215 -0.085 1.295 0.255 ;
        RECT 1.295 -0.085 1.780 0.085 ;
        RECT 1.780 -0.085 1.870 0.305 ;
        RECT 1.870 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.445 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.870 0.125 1.225 ;
      RECT 0.125 0.870 0.205 0.950 ;
      RECT 0.205 0.325 0.230 0.950 ;
      RECT 0.230 0.180 0.280 0.950 ;
      RECT 0.205 1.020 0.345 1.225 ;
      RECT 0.280 0.870 0.435 0.950 ;
      RECT 0.280 0.180 0.530 0.390 ;
      RECT 0.435 0.870 0.530 1.075 ;
      RECT 0.345 1.145 0.780 1.225 ;
      RECT 0.780 1.035 0.860 1.225 ;
      RECT 0.595 0.175 1.125 0.245 ;
      RECT 0.530 0.320 1.385 0.390 ;
      RECT 1.385 0.155 1.440 0.390 ;
      RECT 1.440 0.155 1.520 0.675 ;
      RECT 0.860 1.035 1.520 1.115 ;
      RECT 1.585 0.190 1.610 0.325 ;
      RECT 1.050 0.825 1.610 0.915 ;
      RECT 1.610 0.190 1.690 0.915 ;
  END
END SACELEM1X4

MACRO SACELEM2X2
  CLASS CORE ;
  FOREIGN SACELEM2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.660 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER metal1 ;
        RECT 0.210 0.750 0.560 0.885 ;
        RECT 0.560 0.750 0.755 0.955 ;
        RECT 0.755 0.875 1.420 0.955 ;
    END
  END A
  PIN M1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 1.700 0.455 2.030 0.665 ;
    END
  END M1
  PIN M2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025250 ;
    PORT
      LAYER metal1 ;
        RECT 1.510 0.735 1.720 0.945 ;
    END
  END M2
  PIN P1
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.027250 ;
    PORT
      LAYER metal1 ;
        RECT 0.560 0.455 0.770 0.665 ;
    END
  END P1
  PIN P2
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.027250 ;
    PORT
      LAYER metal1 ;
        RECT 0.180 0.455 0.470 0.660 ;
    END
  END P2
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.081400 ;
    PORT
      LAYER metal1 ;
        RECT 2.325 0.780 2.525 0.875 ;
        RECT 2.525 0.150 2.615 1.155 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052500 ;
    PORT
      LAYER metal1 ;
        RECT 0.860 0.480 0.965 0.805 ;
        RECT 0.965 0.595 1.150 0.805 ;
        RECT 1.150 0.595 1.380 0.685 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.820 1.485 ;
        RECT 0.820 1.180 1.000 1.485 ;
        RECT 1.000 1.315 2.325 1.485 ;
        RECT 2.325 0.965 2.420 1.485 ;
        RECT 2.420 1.315 2.660 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 1.090 0.085 ;
        RECT 1.090 -0.085 1.380 0.195 ;
        RECT 1.380 -0.085 1.880 0.085 ;
        RECT 1.880 -0.085 2.015 0.195 ;
        RECT 2.015 -0.085 2.325 0.085 ;
        RECT 2.325 -0.085 2.420 0.485 ;
        RECT 2.420 -0.085 2.660 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.310 0.115 1.050 ;
      RECT 0.115 0.970 0.125 1.050 ;
      RECT 0.125 0.970 0.345 1.210 ;
      RECT 0.065 0.175 1.000 0.245 ;
      RECT 0.115 0.310 1.420 0.390 ;
      RECT 1.055 0.455 1.510 0.530 ;
      RECT 1.510 0.285 1.610 0.530 ;
      RECT 1.285 1.155 1.820 1.225 ;
      RECT 0.345 1.020 1.910 1.090 ;
      RECT 1.910 1.020 1.920 1.225 ;
      RECT 1.920 0.740 2.055 1.225 ;
      RECT 1.610 0.285 2.145 0.365 ;
      RECT 2.145 0.285 2.235 1.240 ;
  END
END SACELEM2X2

MACRO SNCL2W11OF2X1
  CLASS CORE ;
  FOREIGN SNCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.130 0.740 0.265 0.955 ;
        RECT 0.265 0.875 1.340 0.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.320 0.585 0.995 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 1.955 0.245 2.045 0.945 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049000 ;
    PORT
      LAYER metal1 ;
        RECT 0.520 0.730 1.085 0.810 ;
        RECT 1.085 0.585 1.165 0.810 ;
        RECT 1.165 0.585 1.410 0.720 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.240 1.485 ;
        RECT 0.240 1.225 0.375 1.485 ;
        RECT 0.375 1.315 1.400 1.485 ;
        RECT 1.400 1.225 1.675 1.485 ;
        RECT 1.675 1.315 1.785 1.485 ;
        RECT 1.785 0.670 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.055 0.085 ;
        RECT 0.055 -0.085 0.145 0.195 ;
        RECT 0.145 -0.085 0.435 0.085 ;
        RECT 0.435 -0.085 0.525 0.195 ;
        RECT 0.525 -0.085 1.165 0.085 ;
        RECT 1.165 -0.085 1.340 0.160 ;
        RECT 1.340 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.865 0.495 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.240 0.175 0.345 0.365 ;
      RECT 0.045 1.045 0.610 1.135 ;
      RECT 0.345 0.285 0.615 0.365 ;
      RECT 0.615 0.175 0.705 0.365 ;
      RECT 0.820 0.175 0.955 0.330 ;
      RECT 0.955 0.250 1.430 0.330 ;
      RECT 0.785 0.415 1.475 0.495 ;
      RECT 1.475 0.415 1.555 0.945 ;
      RECT 1.430 0.175 1.620 0.330 ;
      RECT 0.820 1.045 1.620 1.135 ;
      RECT 1.620 0.175 1.695 1.135 ;
  END
END SNCL2W11OF2X1

MACRO SNCL2W11OF2X2
  CLASS CORE ;
  FOREIGN SNCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.090 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.205 0.680 0.310 0.955 ;
        RECT 0.310 0.875 0.625 0.955 ;
        RECT 0.625 0.875 0.705 1.180 ;
        RECT 0.705 0.875 1.225 0.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.290 0.385 0.400 0.590 ;
        RECT 0.400 0.385 0.565 0.665 ;
        RECT 0.565 0.580 1.035 0.665 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.079200 ;
    PORT
      LAYER metal1 ;
        RECT 1.955 0.245 2.045 1.080 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.049500 ;
    PORT
      LAYER metal1 ;
        RECT 0.555 0.730 1.130 0.805 ;
        RECT 1.130 0.580 1.415 0.805 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.220 1.485 ;
        RECT 0.220 1.190 0.310 1.485 ;
        RECT 0.310 1.315 1.360 1.485 ;
        RECT 1.360 1.225 1.645 1.485 ;
        RECT 1.645 1.315 1.785 1.485 ;
        RECT 1.785 0.665 1.865 1.485 ;
        RECT 1.865 1.315 2.090 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.195 ;
        RECT 0.130 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.535 0.160 ;
        RECT 0.535 -0.085 1.165 0.085 ;
        RECT 1.165 -0.085 1.310 0.160 ;
        RECT 1.310 -0.085 1.785 0.085 ;
        RECT 1.785 -0.085 1.865 0.490 ;
        RECT 1.865 -0.085 2.090 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.045 0.920 0.125 1.235 ;
      RECT 0.125 1.020 0.130 1.235 ;
      RECT 0.220 0.175 0.310 0.320 ;
      RECT 0.130 1.020 0.400 1.100 ;
      RECT 0.400 1.020 0.535 1.225 ;
      RECT 0.310 0.250 0.625 0.320 ;
      RECT 0.625 0.175 0.735 0.320 ;
      RECT 0.825 0.175 0.925 0.330 ;
      RECT 0.925 0.250 1.400 0.330 ;
      RECT 0.685 0.410 1.480 0.490 ;
      RECT 1.480 0.410 1.560 0.940 ;
      RECT 1.400 0.175 1.625 0.330 ;
      RECT 0.790 1.045 1.625 1.135 ;
      RECT 1.625 0.175 1.695 1.135 ;
  END
END SNCL2W11OF2X2

MACRO SNCL2W11OF2X4
  CLASS CORE ;
  FOREIGN SNCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.058500 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.665 0.390 0.945 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.058500 ;
    PORT
      LAYER metal1 ;
        RECT 0.120 0.505 0.560 0.585 ;
        RECT 0.560 0.505 0.895 0.805 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.102950 ;
    PORT
      LAYER metal1 ;
        RECT 1.960 0.230 2.055 1.120 ;
    END
  END Q
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.028250 ;
    PORT
      LAYER metal1 ;
        RECT 1.130 0.725 1.340 0.945 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.125 1.485 ;
        RECT 0.125 1.315 0.440 1.485 ;
        RECT 0.440 1.190 0.530 1.485 ;
        RECT 0.530 1.315 1.780 1.485 ;
        RECT 1.780 0.705 1.870 1.485 ;
        RECT 1.870 1.315 2.145 1.485 ;
        RECT 2.145 0.705 2.235 1.485 ;
        RECT 2.235 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.385 ;
        RECT 0.125 -0.085 0.440 0.085 ;
        RECT 0.440 -0.085 0.530 0.245 ;
        RECT 0.530 -0.085 1.380 0.085 ;
        RECT 1.380 -0.085 1.515 0.360 ;
        RECT 1.515 -0.085 1.780 0.085 ;
        RECT 1.780 -0.085 1.870 0.305 ;
        RECT 1.870 -0.085 2.145 0.085 ;
        RECT 2.145 -0.085 2.235 0.520 ;
        RECT 2.235 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.215 0.175 0.350 0.415 ;
      RECT 0.215 1.020 0.350 1.225 ;
      RECT 0.350 0.335 0.620 0.415 ;
      RECT 0.350 1.020 0.620 1.100 ;
      RECT 0.620 0.175 0.700 0.415 ;
      RECT 0.620 1.020 0.700 1.225 ;
      RECT 0.790 0.895 0.895 1.080 ;
      RECT 0.790 0.315 1.005 0.415 ;
      RECT 0.700 0.175 1.085 0.250 ;
      RECT 1.005 0.315 1.085 0.660 ;
      RECT 0.700 1.145 1.085 1.225 ;
      RECT 0.895 1.010 1.185 1.080 ;
      RECT 1.085 0.315 1.280 0.385 ;
      RECT 1.185 1.010 1.320 1.225 ;
      RECT 1.085 0.585 1.430 0.660 ;
      RECT 1.430 0.585 1.520 1.225 ;
      RECT 1.150 0.450 1.585 0.520 ;
      RECT 1.585 0.230 1.610 0.520 ;
      RECT 1.585 0.690 1.610 0.980 ;
      RECT 1.610 0.230 1.690 0.980 ;
  END
END SNCL2W11OF2X4

MACRO SRNCL2W11OF2X1
  CLASS CORE ;
  FOREIGN SRNCL2W11OF2X1 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.510 0.760 ;
        RECT 0.510 0.525 0.600 0.615 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.115 0.855 0.690 0.945 ;
        RECT 0.690 0.600 0.815 0.945 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.039600 ;
    PORT
      LAYER metal1 ;
        RECT 2.150 0.525 2.335 0.655 ;
        RECT 2.335 0.355 2.425 1.020 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 0.915 0.665 1.270 0.945 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 1.360 0.665 1.650 1.020 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.035 0.130 1.485 ;
        RECT 0.130 1.315 0.445 1.485 ;
        RECT 0.445 1.180 0.535 1.485 ;
        RECT 0.535 1.315 1.085 1.485 ;
        RECT 1.085 1.290 1.285 1.485 ;
        RECT 1.285 1.315 2.150 1.485 ;
        RECT 2.150 0.745 2.240 1.485 ;
        RECT 2.240 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.420 ;
        RECT 0.130 -0.085 0.445 0.085 ;
        RECT 0.445 -0.085 0.535 0.280 ;
        RECT 0.535 -0.085 1.780 0.085 ;
        RECT 1.780 -0.085 1.915 0.275 ;
        RECT 1.915 -0.085 2.150 0.085 ;
        RECT 2.150 -0.085 2.240 0.435 ;
        RECT 2.240 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.180 0.355 0.435 ;
      RECT 0.220 1.020 0.355 1.225 ;
      RECT 0.355 0.355 0.915 0.435 ;
      RECT 0.915 0.320 1.130 0.435 ;
      RECT 0.355 1.020 1.130 1.090 ;
      RECT 0.725 0.175 1.195 0.255 ;
      RECT 1.195 0.175 1.275 0.450 ;
      RECT 0.970 0.525 1.340 0.595 ;
      RECT 1.340 0.175 1.420 0.595 ;
      RECT 0.725 1.155 1.510 1.225 ;
      RECT 1.485 0.315 1.565 0.600 ;
      RECT 1.420 0.175 1.630 0.250 ;
      RECT 1.630 0.175 1.710 0.445 ;
      RECT 1.565 0.520 1.740 0.600 ;
      RECT 1.600 1.110 1.740 1.200 ;
      RECT 1.740 0.520 1.820 1.200 ;
      RECT 1.820 0.520 1.880 0.725 ;
      RECT 1.710 0.365 1.970 0.445 ;
      RECT 1.970 0.365 2.060 1.020 ;
  END
END SRNCL2W11OF2X1

MACRO SRNCL2W11OF2X2
  CLASS CORE ;
  FOREIGN SRNCL2W11OF2X2 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.280 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.510 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.125 0.825 0.600 0.905 ;
        RECT 0.600 0.525 0.890 0.905 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.076650 ;
    PORT
      LAYER metal1 ;
        RECT 2.010 0.640 2.150 0.875 ;
        RECT 2.150 0.245 2.155 0.875 ;
        RECT 2.155 0.245 2.235 1.170 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 1.010 0.525 1.300 0.735 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.026000 ;
    PORT
      LAYER metal1 ;
        RECT 1.390 0.525 1.650 0.735 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.030 0.125 1.485 ;
        RECT 0.125 1.315 0.400 1.485 ;
        RECT 0.400 1.185 0.535 1.485 ;
        RECT 0.535 1.315 1.080 1.485 ;
        RECT 1.080 1.290 1.270 1.485 ;
        RECT 1.270 1.315 1.985 1.485 ;
        RECT 1.985 0.965 2.065 1.485 ;
        RECT 2.065 1.315 2.280 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.130 0.435 ;
        RECT 0.130 -0.085 0.400 0.085 ;
        RECT 0.400 -0.085 0.535 0.260 ;
        RECT 0.535 -0.085 1.585 0.085 ;
        RECT 1.585 -0.085 1.665 0.275 ;
        RECT 1.665 -0.085 1.985 0.085 ;
        RECT 1.985 -0.085 2.065 0.305 ;
        RECT 2.065 -0.085 2.280 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.220 0.160 0.310 0.435 ;
      RECT 0.205 0.985 0.310 1.225 ;
      RECT 0.310 0.355 0.900 0.435 ;
      RECT 0.900 0.335 1.115 0.435 ;
      RECT 0.310 0.985 1.115 1.065 ;
      RECT 0.700 0.175 1.270 0.260 ;
      RECT 0.700 1.130 1.330 1.210 ;
      RECT 1.330 1.000 1.460 1.210 ;
      RECT 1.360 0.175 1.495 0.435 ;
      RECT 0.985 0.825 1.545 0.905 ;
      RECT 1.545 0.825 1.625 1.205 ;
      RECT 1.495 0.355 1.715 0.435 ;
      RECT 1.715 0.355 1.785 0.910 ;
      RECT 1.755 0.175 1.850 0.265 ;
      RECT 1.625 1.000 1.850 1.205 ;
      RECT 1.850 0.175 1.920 1.205 ;
  END
END SRNCL2W11OF2X2

MACRO SRNCL2W11OF2X4
  CLASS CORE ;
  FOREIGN SRNCL2W11OF2X4 0.000 0.000 ;
  ORIGIN 0.000 0.000 ;
  SYMMETRY X Y ;
  SITE core10T ;
  SIZE 2.470 BY 1.400 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.440 0.485 0.920 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.052000 ;
    PORT
      LAYER metal1 ;
        RECT 0.060 0.525 0.350 0.905 ;
        RECT 0.350 0.825 0.830 0.905 ;
    END
  END B
  PIN Q
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.105850 ;
    PORT
      LAYER metal1 ;
        RECT 2.140 0.245 2.230 1.235 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025000 ;
    PORT
      LAYER metal1 ;
        RECT 1.120 0.455 1.530 0.665 ;
    END
  END RN
  PIN S
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.025500 ;
    PORT
      LAYER metal1 ;
        RECT 1.320 0.735 1.555 0.945 ;
    END
  END S
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 1.315 0.045 1.485 ;
        RECT 0.045 1.025 0.125 1.485 ;
        RECT 0.125 1.315 0.435 1.485 ;
        RECT 0.435 1.165 0.525 1.485 ;
        RECT 0.525 1.315 1.070 1.485 ;
        RECT 1.070 1.290 1.260 1.485 ;
        RECT 1.260 1.315 1.960 1.485 ;
        RECT 1.960 1.170 2.050 1.485 ;
        RECT 2.050 1.315 2.335 1.485 ;
        RECT 2.335 0.830 2.425 1.485 ;
        RECT 2.425 1.315 2.470 1.485 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.000 -0.085 0.045 0.085 ;
        RECT 0.045 -0.085 0.125 0.420 ;
        RECT 0.125 -0.085 0.415 0.085 ;
        RECT 0.415 -0.085 0.550 0.245 ;
        RECT 0.550 -0.085 1.545 0.085 ;
        RECT 1.545 -0.085 1.765 0.195 ;
        RECT 1.765 -0.085 1.960 0.085 ;
        RECT 1.960 -0.085 2.050 0.470 ;
        RECT 2.050 -0.085 2.335 0.085 ;
        RECT 2.335 -0.085 2.425 0.460 ;
        RECT 2.425 -0.085 2.470 0.085 ;
    END
  END VSS
  OBS
    LAYER metal1 ;
      RECT 0.210 0.995 0.345 1.225 ;
      RECT 0.215 0.180 0.350 0.390 ;
      RECT 0.345 0.995 1.105 1.075 ;
      RECT 0.350 0.320 1.120 0.390 ;
      RECT 1.010 0.770 1.170 0.905 ;
      RECT 1.170 0.770 1.250 1.080 ;
      RECT 0.730 0.175 1.275 0.255 ;
      RECT 1.365 0.175 1.455 0.365 ;
      RECT 0.705 1.145 1.480 1.225 ;
      RECT 1.250 1.010 1.545 1.080 ;
      RECT 1.545 1.010 1.595 1.195 ;
      RECT 1.455 0.285 1.645 0.365 ;
      RECT 1.645 0.285 1.715 0.965 ;
      RECT 1.715 0.730 1.780 0.965 ;
      RECT 1.780 0.400 1.870 0.640 ;
      RECT 1.780 0.730 1.870 0.865 ;
      RECT 1.595 1.030 1.870 1.195 ;
      RECT 1.870 0.560 1.960 0.640 ;
      RECT 1.870 1.030 1.960 1.105 ;
      RECT 1.960 0.560 2.050 1.105 ;
  END
END SRNCL2W11OF2X4

END LIBRARY
##############################################################################
#                                                                            #
# End of file.                                                               #
#                                                                            #
##############################################################################

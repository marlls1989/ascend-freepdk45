.SUBCKT ACELEM1X1 A M P Q VDD VSS
*.PININFO A:I M:I P:I Q:O VDD:P VSS:G
M_i_0 net_6 M VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_1 VSS A net_6 VSS NMOS_VTL W=180n L=50n M=1
M_i_2 net_6 net_8 net_7 VSS NMOS_VTL W=180n L=50n M=1
M_i_3 net_7 A net_10 VSS NMOS_VTL W=180n L=50n M=1
M_i_4 net_10 P VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_5 net_8 net_7 VSS VSS NMOS_VTL W=155n L=50n M=1
M_i_6 VSS net_7 Q VSS NMOS_VTL W=155n L=50n M=1
M_i_7 VDD M net_11 VDD PMOS_VTL W=240n L=50n M=1
M_i_8 net_11 A net_7 VDD PMOS_VTL W=240n L=50n M=1
M_i_9 net_7 net_8 net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_10 net_9 A VDD VDD PMOS_VTL W=240n L=50n M=1
M_i_11 VDD P net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_12 net_8 net_7 VDD VDD PMOS_VTL W=215n L=50n M=1
M_i_13 VDD net_7 Q VDD PMOS_VTL W=215n L=50n M=1
.ENDS
.SUBCKT ACELEM1X2 A M P Q VDD VSS
*.PININFO A:I M:I P:I Q:O VDD:P VSS:G
M_i_0 net_6 M VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_1 VSS A net_6 VSS NMOS_VTL W=180n L=50n M=1
M_i_2 net_6 net_8 net_7 VSS NMOS_VTL W=180n L=50n M=1
M_i_3 net_7 A net_10 VSS NMOS_VTL W=180n L=50n M=1
M_i_4 net_10 P VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_5 net_8 net_7 VSS VSS NMOS_VTL W=155n L=50n M=1
M_i_6 VSS net_7 Q VSS NMOS_VTL W=305n L=50n M=1
M_i_7 VDD M net_11 VDD PMOS_VTL W=240n L=50n M=1
M_i_8 net_11 A net_7 VDD PMOS_VTL W=240n L=50n M=1
M_i_9 net_7 net_8 net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_10 net_9 A VDD VDD PMOS_VTL W=240n L=50n M=1
M_i_11 VDD P net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_12 net_8 net_7 VDD VDD PMOS_VTL W=215n L=50n M=1
M_i_13 VDD net_7 Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT ACELEM1X4 A M P Q VDD VSS
*.PININFO A:I M:I P:I Q:O VDD:P VSS:G
M_i_0 net_6 M VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_1 VSS A net_6 VSS NMOS_VTL W=180n L=50n M=1
M_i_2 net_6 net_8 net_7 VSS NMOS_VTL W=180n L=50n M=1
M_i_3 net_7 A net_10 VSS NMOS_VTL W=180n L=50n M=1
M_i_4 net_10 P VSS VSS NMOS_VTL W=180n L=50n M=1
M_i_5 net_8 net_7 VSS VSS NMOS_VTL W=155n L=50n M=1
M_i_6 VSS net_7 Q VSS NMOS_VTL W=305n L=50n M=1
M_i_7 VSS net_7 Q VSS NMOS_VTL W=305n L=50n M=1
M_i_8 VDD M net_11 VDD PMOS_VTL W=240n L=50n M=1
M_i_9 net_11 A net_7 VDD PMOS_VTL W=240n L=50n M=1
M_i_10 net_7 net_8 net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_11 net_9 A VDD VDD PMOS_VTL W=240n L=50n M=1
M_i_12 VDD P net_9 VDD PMOS_VTL W=240n L=50n M=1
M_i_13 net_8 net_7 VDD VDD PMOS_VTL W=215n L=50n M=1
M_i_14 VDD net_7 Q VDD PMOS_VTL W=415n L=50n M=1
M_i_15 VDD net_7 Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT FILL1 VDD VSS
*.PININFO VDD:P VSS:G
.ENDS
.SUBCKT FILLTIE VDD VSS
*.PININFO VDD:P VSS:G
.ENDS
.SUBCKT INCL1W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D Q VDD PMOS_VTL W=340n L=50n M=1
MNI0 Q A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI1 Q B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 Q C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 Q D VSS VSS NMOS_VTL W=180n L=50n M=1
.ENDS
.SUBCKT INCL1W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C Q VDD PMOS_VTL W=305n L=50n M=1
MNI0 Q A VSS VSS NMOS_VTL W=115n L=50n M=1
MNI1 Q B VSS VSS NMOS_VTL W=115n L=50n M=1
MNI2 Q C VSS VSS NMOS_VTL W=115n L=50n M=1
.ENDS
.SUBCKT INCL1W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 Q B VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_0 VSS A Q VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 net_0 B VDD VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_2 Q A net_0 VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
.ENDS
.SUBCKT INCL1W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 Q B VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_0 VSS A Q VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 net_0 B VDD VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_2 Q A net_0 VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
.ENDS
.SUBCKT INCL1W1OF1X1 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPO0 VDD A Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q A VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCL1W1OF1X2 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPO0 VDD A Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q A VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL1W1OF1X4 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPO0 VDD A Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD A Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q A VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q A VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL2W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT INCL2W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL2W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL2W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCL2W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL2W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL3W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCL3W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL3W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL3W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT INCL3W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL3W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCL4W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCL4W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL4W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP1W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 Q A VDD VDD PMOS_VTL W=250n L=50n M=1
MPI1 Q B VDD VDD PMOS_VTL W=250n L=50n M=1
MPI2 Q C VDD VDD PMOS_VTL W=250n L=50n M=1
MPI3 Q D VDD VDD PMOS_VTL W=250n L=50n M=1
MNI0 Q D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
.ENDS
.SUBCKT INCLP1W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A Q VDD PMOS_VTL W=205n L=50n M=1
MPI1 VDD B Q VDD PMOS_VTL W=205n L=50n M=1
MPI2 VDD C Q VDD PMOS_VTL W=205n L=50n M=1
MNI0 Q C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT INCLP1W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 net_0 B VSS VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_0 Q A net_0 VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_3 Q B VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_2 VDD A Q VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
.ENDS
.SUBCKT INCLP1W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 net_0 B VSS VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_0 Q A net_0 VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_3 Q B VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
M_i_2 VDD A Q VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
.ENDS
.SUBCKT INCLP2W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT INCLP2W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCLP2W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCLP2W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCLP2W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP2W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP3W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCLP3W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCLP3W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT INCLP4W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCLP4W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP4W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 PREQ D VSS VSS NMOS_VTL W=180n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL1W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 PREQ D VSS VSS NMOS_VTL W=180n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=115n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=115n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=115n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL1W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=115n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=115n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=115n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=115n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=115n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=115n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 Q_neg B VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_0 VSS A Q_neg VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 net_0 B VDD VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_2 Q_neg A net_0 VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_4 Q Q_neg VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 Q Q_neg VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
.ENDS
.SUBCKT NCL1W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_1 Q_neg B VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_0 VSS A Q_neg VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 net_0 B VDD VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_2 Q_neg A net_0 VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_4 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
.ENDS
.SUBCKT NCL1W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_0 Q_neg B VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_1 VSS A Q_neg VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_2 net_0 B VDD VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_3 Q_neg A net_0 VDD PMOS_VTL W=250n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_4 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_6 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_7 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
.ENDS
.SUBCKT NCL1W1OF1X1 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL1W1OF1X2 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W1OF1X4 A Q VDD VSS
*.PININFO A:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL2W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT NCL2W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL2W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL2W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL2W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL2W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 C PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL3W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT NCL3W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL3W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL3W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT NCL3W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL3W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD C pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ A nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCL3W3111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL3W3111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL4W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCL4W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL4W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLAO22OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLAO22OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLAO22OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 B ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLOA22OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph02 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLOA22OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph02 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLOA22OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph02 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP1W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 PREQ A VDD VDD PMOS_VTL W=250n L=50n M=1
MPI1 PREQ B VDD VDD PMOS_VTL W=250n L=50n M=1
MPI2 PREQ C VDD VDD PMOS_VTL W=250n L=50n M=1
MPI3 PREQ D VDD VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP1W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 PREQ A VDD VDD PMOS_VTL W=250n L=50n M=1
MPI1 PREQ B VDD VDD PMOS_VTL W=250n L=50n M=1
MPI2 PREQ C VDD VDD PMOS_VTL W=250n L=50n M=1
MPI3 PREQ D VDD VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP1W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 PREQ A VDD VDD PMOS_VTL W=250n L=50n M=1
MPI1 PREQ B VDD VDD PMOS_VTL W=250n L=50n M=1
MPI2 PREQ C VDD VDD PMOS_VTL W=250n L=50n M=1
MPI3 PREQ D VDD VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP1W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI1 VDD B PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI2 VDD C PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP1W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI1 VDD B PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI2 VDD C PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP1W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI1 VDD B PREQ VDD PMOS_VTL W=205n L=50n M=1
MPI2 VDD C PREQ VDD PMOS_VTL W=205n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP1W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_2 net_0 A Q_neg VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_3 VSS B net_0 VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_0 Q Q_neg VSS VSS NMOS_VTL W=155n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_4 Q_neg A VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 VDD B Q_neg VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_1 Q Q_neg VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
.ENDS
.SUBCKT NCLP1W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_2 net_0 A Q_neg VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_3 VSS B net_0 VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_0 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_4 Q_neg A VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 VDD B Q_neg VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_1 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
.ENDS
.SUBCKT NCLP1W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_0 net_0 A Q_neg VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_1 VSS B net_0 VSS NMOS_VTL W=180n L=50n M=1 AD=0.016200P AS=0.016200P PD=0.360000U PS=0.360000U
M_i_2 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 Q Q_neg VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_4 Q_neg A VDD VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_5 VDD B Q_neg VDD PMOS_VTL W=205n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_6 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
M_i_7 Q Q_neg VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.021012P AS=0.021012P PD=0.410000U PS=0.410000U
.ENDS
.SUBCKT NCLP2W11OF2X1 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT NCLP2W11OF2X2 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCLP2W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCLP2W211OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP2W211OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP2W211OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD B pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS C nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ A NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP3W111OF3X1 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT NCLP3W111OF3X2 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCLP3W111OF3X4 A B C Q VDD VSS
*.PININFO A:I B:I C:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI2 pl01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ C nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 B nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT NCLP4W1111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP4W1111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP4W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP4W3111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP4W3111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLPAO22OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH3 nh01 C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh01 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLPAO22OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH3 nh01 C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh01 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLPOA22OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD B pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 nh01 B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh02 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh02 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLPOA22OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD B pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 nh01 B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh02 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh02 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLPOA22OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD B pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 nh01 B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh02 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh02 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT PULLDOWN Q VDD VSS
*.PININFO VDD:P VSS:G
M_i_0 VSS Q Q VSS NMOS_VTL W=295n L=50n M=1
.ENDS
.SUBCKT PULLUP Q VDD VSS
*.PININFO VDD:P VSS:G
M_i_0 VDD Q Q VDD PMOS_VTL W=405n L=50n M=1
.ENDS
.SUBCKT RACELEM1X1 A M P RN Q VDD VSS
*.PININFO A:I M:I P:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI1 VDD P pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A NNET VSS NMOS_VTL W=205n L=50n M=1
MNG0 NNET RN PREQ VSS NMOS_VTL W=205n L=50n M=1
MPH0 NNET IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT RACELEM1X2 A M P RN Q VDD VSS
*.PININFO A:I M:I P:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI1 VDD P pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A NNET VSS NMOS_VTL W=205n L=50n M=1
MNG0 NNET RN PREQ VSS NMOS_VTL W=205n L=50n M=1
MPH0 NNET IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT RACELEM1X4 A M P RN Q VDD VSS
*.PININFO A:I M:I P:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI1 VDD P pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A NNET VSS NMOS_VTL W=205n L=50n M=1
MNG0 NNET RN PREQ VSS NMOS_VTL W=205n L=50n M=1
MPH0 NNET IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT RACELEM2X1 A M1 M2 P1 P2 RN Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD P1 pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 P2 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 RN PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M1 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 M2 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 RN nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 PREQ P1 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 PREQ P2 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH4 PREQ A nh01 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=115n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT RACELEM2X2 A M1 M2 P1 P2 RN Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD P1 pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 P2 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 RN PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M1 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 M2 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 RN nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 PREQ P1 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 PREQ P2 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH4 PREQ A nh01 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT RACELEM2X4 A M1 M2 P1 P2 RN Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I RN:I Q:O VDD:P VSS:G
MPI0 VDD RN PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI1 VDD P1 pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl00 P2 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 RN PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 M1 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 M2 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 RN nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 PREQ P1 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 PREQ P2 nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH4 PREQ A nh01 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT RNCL2W11OF2X1 A B RN Q VDD VSS
*.PININFO A:I B:I RN:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT RNCL2W11OF2X2 A B RN Q VDD VSS
*.PININFO A:I B:I RN:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT RNCL2W11OF2X4 A B RN Q VDD VSS
*.PININFO A:I B:I RN:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT RSNCL2W11OF2X1 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 NNET S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT RSNCL2W11OF2X2 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 NNET S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT RSNCL2W11OF2X4 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 NNET S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SACELEM1X1 A M P S Q VDD VSS
*.PININFO A:I M:I P:I S:I Q:O VDD:P VSS:G
MPI0 VDD P pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 A PNET VDD PMOS_VTL W=305n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A PREQ VSS NMOS_VTL W=180n L=50n M=1
MNI2 VSS S PREQ VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT SACELEM1X2 A M P S Q VDD VSS
*.PININFO A:I M:I P:I S:I Q:O VDD:P VSS:G
MPI0 VDD P pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 A PNET VDD PMOS_VTL W=305n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A PREQ VSS NMOS_VTL W=180n L=50n M=1
MNI2 VSS S PREQ VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT SACELEM1X4 A M P S Q VDD VSS
*.PININFO A:I M:I P:I S:I Q:O VDD:P VSS:G
MPI0 VDD P pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 A PNET VDD PMOS_VTL W=305n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 VSS M nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A PREQ VSS NMOS_VTL W=180n L=50n M=1
MNI2 VSS S PREQ VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 M VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS P nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
.ENDS
.SUBCKT SACELEM2X2 A M1 M2 P1 P2 S Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I S:I Q:O VDD:P VSS:G
MPI0 VDD S pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 P1 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 P2 pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A PREQ VSS NMOS_VTL W=235n L=50n M=1
MNI3 VSS S PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 S ph01 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph01 M1 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph01 M2 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph01 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=205n L=50n M=1
MNH1 PREQ S nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 PREQ P1 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 PREQ P2 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH4 PREQ A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SNCL2W11OF2X1 A B S Q VDD VSS
*.PININFO A:I B:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT SNCL2W11OF2X2 A B S Q VDD VSS
*.PININFO A:I B:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SNCL2W11OF2X4 A B S Q VDD VSS
*.PININFO A:I B:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ B nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SRNCL2W11OF2X1 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT SRNCL2W11OF2X2 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SRNCL2W11OF2X4 A B RN S Q VDD VSS
*.PININFO A:I B:I RN:I S:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B PNET VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD RN PNET VDD PMOS_VTL W=305n L=50n M=1
MNI0 NNET B nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 A VSS VSS NMOS_VTL W=205n L=50n M=1
MNI2 PREQ S VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PNET IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph00 A VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph00 B VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ NNET VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPG0 PNET S PREQ VDD PMOS_VTL W=305n L=50n M=1
MNG0 PREQ RN NNET VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL1W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_0 Q B VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_1 Q B VSS VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_2 VSS A Q VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_3 VSS A Q VSS NMOS_VTL W=305n L=50n M=1 AD=0.012013P AS=0.012013P PD=0.310000U PS=0.310000U
M_i_4 net_0 B VDD VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_5 net_1 B VDD VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_6 Q A net_0 VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
M_i_7 Q A net_1 VDD PMOS_VTL W=500n L=50n M=1 AD=0.031250P AS=0.031250P PD=0.500000U PS=0.500000U
.ENDS
.SUBCKT INCL3W2211OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=115n L=50n M=1
.ENDS
.SUBCKT INCL3W2211OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL3W2211OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL3W3111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCL3W3111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCL3W3111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B VDD VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C VDD VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D VDD VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP1W11OF2X4 A B Q VDD VSS
*.PININFO A:I B:I Q:O VDD:P VSS:G
M_i_0 net_0 B VSS VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_1 net_1 B VSS VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_2 Q A net_0 VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_3 Q A net_1 VSS NMOS_VTL W=360n L=50n M=1 AD=0.064800P AS=0.064800P PD=0.720000U PS=0.720000U
M_i_4 Q B VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
M_i_5 Q B VDD VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
M_i_6 VDD A Q VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
M_i_7 VDD A Q VDD PMOS_VTL W=415n L=50n M=1 AD=0.086113P AS=0.086113P PD=0.830000U PS=0.830000U
.ENDS
.SUBCKT INCLP4W2211OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCLP4W2211OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP4W2211OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP4W3111OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT INCLP4W3111OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT INCLP4W3111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD IQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q IQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL1W1111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI2 PREQ C VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 PREQ D VSS VSS NMOS_VTL W=180n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL3W2211OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=115n L=50n M=1
.ENDS
.SUBCKT NCL3W2211OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL3W2211OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 PREQ C nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl00 B VSS VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl00 A VSS VSS NMOS_VTL W=180n L=50n M=1
MNI4 PREQ B nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI5 nl01 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=340n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=340n L=50n M=1
MPH2 ph01 B ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH3 ph00 C ph02 VDD PMOS_VTL W=340n L=50n M=1
MPH4 ph02 D ph03 VDD PMOS_VTL W=340n L=50n M=1
MPH5 ph03 A VDD VDD PMOS_VTL W=340n L=50n M=1
MPH6 ph03 B VDD VDD PMOS_VTL W=340n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=180n L=50n M=1
MNH1 VSS A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 VSS B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 VSS C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 VSS D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCL3W3111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 C pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=205n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=205n L=50n M=1
MNI2 nl01 B VSS VSS NMOS_VTL W=205n L=50n M=1
MNI3 PREQ A VSS VSS NMOS_VTL W=205n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=305n L=50n M=1
MPH1 ph00 A ph01 VDD PMOS_VTL W=305n L=50n M=1
MPH2 ph01 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH3 ph01 C PREQ VDD PMOS_VTL W=305n L=50n M=1
MPH4 ph01 D PREQ VDD PMOS_VTL W=305n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH3 PREQ C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 PREQ D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP4W2211OF4X1 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
.ENDS
.SUBCKT NCLP4W2211OF4X2 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP4W2211OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=305n L=50n M=1
MPI1 pl00 B pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=305n L=50n M=1
MPI3 pl01 D pl03 VDD PMOS_VTL W=305n L=50n M=1
MPI4 pl03 A PREQ VDD PMOS_VTL W=305n L=50n M=1
MPI5 pl03 B PREQ VDD PMOS_VTL W=305n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=180n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=180n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=180n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=180n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A VDD VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 nh01 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS B nh01 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS C nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS D nh02 VSS NMOS_VTL W=205n L=50n M=1
MNH5 nh02 A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH6 nh02 B nh00 VSS NMOS_VTL W=205n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLP4W3111OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=250n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI2 pl00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPI3 pl00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=235n L=50n M=1
MNH1 PREQ A nh00 VSS NMOS_VTL W=235n L=50n M=1
MNH2 PREQ D nh01 VSS NMOS_VTL W=235n L=50n M=1
MNH3 nh01 C nh02 VSS NMOS_VTL W=235n L=50n M=1
MNH4 nh02 B nh00 VSS NMOS_VTL W=235n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT NCLPAO22OF4X4 A B C D Q VDD VSS
*.PININFO A:I B:I C:I D:I Q:O VDD:P VSS:G
MPI0 VDD A pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 B PREQ VDD PMOS_VTL W=340n L=50n M=1
MPI2 VDD C pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl01 D PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 PREQ D nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 C nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 B nl02 VSS NMOS_VTL W=235n L=50n M=1
MNI3 nl02 A VSS VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph00 B PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph00 C PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph00 D PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=180n L=50n M=1
MNH1 PREQ A nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH2 PREQ B nh01 VSS NMOS_VTL W=180n L=50n M=1
MNH3 nh01 C nh00 VSS NMOS_VTL W=180n L=50n M=1
MNH4 nh01 D nh00 VSS NMOS_VTL W=180n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=415n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=305n L=50n M=1
.ENDS
.SUBCKT SACELEM2X1 A M1 M2 P1 P2 S Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I S:I Q:O VDD:P VSS:G
MPI0 VDD S pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 P1 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 P2 pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A PREQ VSS NMOS_VTL W=235n L=50n M=1
MNI3 VSS S PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 PREQ IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 S ph01 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph01 M1 VDD VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph01 M2 VDD VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph01 A VDD VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ PREQ VSS NMOS_VTL W=205n L=50n M=1
MNH1 VSS S nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 VSS P1 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 VSS P2 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH4 VSS A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=205n L=50n M=1
.ENDS
.SUBCKT SACELEM2X4 A M1 M2 P1 P2 S Q VDD VSS
*.PININFO A:I M1:I M2:I P1:I P2:I S:I Q:O VDD:P VSS:G
MPI0 VDD S pl00 VDD PMOS_VTL W=340n L=50n M=1
MPI1 pl00 P1 pl01 VDD PMOS_VTL W=340n L=50n M=1
MPI2 pl01 P2 pl02 VDD PMOS_VTL W=340n L=50n M=1
MPI3 pl02 A PREQ VDD PMOS_VTL W=340n L=50n M=1
MNI0 VSS M1 nl00 VSS NMOS_VTL W=235n L=50n M=1
MNI1 nl00 M2 nl01 VSS NMOS_VTL W=235n L=50n M=1
MNI2 nl01 A PREQ VSS NMOS_VTL W=235n L=50n M=1
MNI3 VSS S PREQ VSS NMOS_VTL W=235n L=50n M=1
MPH0 VDD IQ ph00 VDD PMOS_VTL W=250n L=50n M=1
MPH1 ph00 S ph01 VDD PMOS_VTL W=250n L=50n M=1
MPH2 ph01 M1 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH3 ph01 M2 PREQ VDD PMOS_VTL W=250n L=50n M=1
MPH4 ph01 A PREQ VDD PMOS_VTL W=250n L=50n M=1
MNH0 nh00 IQ VSS VSS NMOS_VTL W=205n L=50n M=1
MNH1 PREQ S nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH2 PREQ P1 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH3 PREQ P2 nh00 VSS NMOS_VTL W=205n L=50n M=1
MNH4 PREQ A nh00 VSS NMOS_VTL W=205n L=50n M=1
MNB0 IQ PREQ VSS VSS NMOS_VTL W=155n L=50n M=1
MPB0 VDD PREQ IQ VDD PMOS_VTL W=205n L=50n M=1
MNO0 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MNO1 Q PREQ VSS VSS NMOS_VTL W=415n L=50n M=1
MPO0 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
MPO1 VDD PREQ Q VDD PMOS_VTL W=305n L=50n M=1
.ENDS
******************************************************************************
*                                                                            *
* End of file.                                                               *
*                                                                            *
******************************************************************************

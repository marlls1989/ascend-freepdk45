
.SUBCKT PULLDOWN Q VDD VSS
*.PININFO VDD:P VSS:G
M_i_0 VSS Q Q VSS NMOS_VTL W=295n L=50n M=1
.ENDS
******************************************************************************
*                                                                            *
* End of file.                                                               *
*                                                                            *
******************************************************************************

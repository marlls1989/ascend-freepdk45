
.SUBCKT PULLUP Q VDD VSS
*.PININFO VDD:P VSS:G
M_i_0 VDD Q Q VDD PMOS_VTL W=405n L=50n M=1
.ENDS
******************************************************************************
*                                                                            *
* End of file.                                                               *
*                                                                            *
******************************************************************************

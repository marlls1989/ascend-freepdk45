
.SUBCKT FILL1 VDD VSS
*.PININFO VDD:P VSS:G
.ENDS
******************************************************************************
*                                                                            *
* End of file.                                                               *
*                                                                            *
******************************************************************************
